library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity vrom is
	port 
	(
		address_a		: in natural range 0 to 8191;
		address_b		: in natural range 0 to 8191;
		clock		: IN STD_LOGIC ;
		q_a		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		q_b		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
end entity;

architecture rtl of vrom is

	-- Build a 2-D array type for the ROM
	-- subtype word_t is std_logic_vector(7 downto 0);
	-- type memory_t is array(8191 downto 0) of word_t;
	subtype word_t is std_logic_vector(0 to 7);
	type memory_t is array(0 to 8191) of word_t;
		
	-- function init_rom
	-- return memory_t is
	-- variable tmp : memory_t := (others => (others => '0'));
	-- begin 
	-- 	for addr_pos in 0 to 8191 loop 
	-- 		-- Initialize each address with the address itself
	-- 		tmp(addr_pos) := std_logic_vector(to_unsigned(addr_pos, 8));
	-- 	end loop;
		
	-- 	return tmp;
	-- end init_rom;
	
	-- Declare the ROM signal and specify a default value. Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	signal rom : memory_t := 
	(
X"03",
X"0f",
X"1f",
X"1f",
X"1c",
X"24",
X"26",
X"66",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"3f",
X"3f",
X"7f",
X"e0",
X"c0",
X"80",
X"fc",
X"80",
X"c0",
X"00",
X"20",
X"00",
X"20",
X"60",
X"00",
X"f0",
X"fc",
X"fe",
X"fe",
X"60",
X"70",
X"18",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"7f",
X"7f",
X"1f",
X"07",
X"00",
X"1e",
X"3f",
X"7f",
X"fc",
X"7c",
X"00",
X"00",
X"e0",
X"f0",
X"f8",
X"f8",
X"fc",
X"fc",
X"f8",
X"c0",
X"c2",
X"67",
X"2f",
X"37",
X"7f",
X"7f",
X"ff",
X"ff",
X"07",
X"07",
X"0f",
X"0f",
X"7f",
X"7e",
X"fc",
X"f0",
X"f8",
X"f8",
X"f0",
X"70",
X"fd",
X"fe",
X"b4",
X"f8",
X"f8",
X"f9",
X"fb",
X"ff",
X"37",
X"36",
X"5c",
X"00",
X"00",
X"01",
X"03",
X"1f",
X"1f",
X"3f",
X"ff",
X"ff",
X"fc",
X"70",
X"70",
X"38",
X"08",
X"24",
X"e3",
X"f0",
X"f8",
X"70",
X"70",
X"38",
X"ff",
X"ff",
X"ff",
X"1f",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"1f",
X"1f",
X"1f",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"07",
X"0f",
X"0f",
X"0e",
X"12",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"1f",
X"00",
X"00",
X"f0",
X"e0",
X"c0",
X"fe",
X"40",
X"60",
X"00",
X"00",
X"00",
X"10",
X"30",
X"00",
X"f8",
X"fe",
X"13",
X"33",
X"30",
X"18",
X"04",
X"0f",
X"1f",
X"1f",
X"1f",
X"3f",
X"3f",
X"1f",
X"07",
X"08",
X"17",
X"17",
X"00",
X"10",
X"7e",
X"3e",
X"00",
X"00",
X"c0",
X"e0",
X"ff",
X"ff",
X"fe",
X"fe",
X"fc",
X"e0",
X"40",
X"a0",
X"3f",
X"3f",
X"3f",
X"1f",
X"1f",
X"1f",
X"1f",
X"1f",
X"37",
X"27",
X"23",
X"03",
X"01",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f0",
X"f8",
X"f8",
X"f8",
X"f8",
X"f8",
X"cc",
X"ff",
X"ff",
X"ff",
X"ff",
X"70",
X"00",
X"08",
X"ff",
X"ff",
X"ff",
X"fe",
X"f0",
X"c0",
X"80",
X"00",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"c0",
X"80",
X"00",
X"fc",
X"fc",
X"f8",
X"78",
X"78",
X"78",
X"7e",
X"7e",
X"10",
X"60",
X"80",
X"00",
X"78",
X"78",
X"7e",
X"7e",
X"00",
X"03",
X"0f",
X"1f",
X"1f",
X"1c",
X"24",
X"26",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"3f",
X"3f",
X"00",
X"e0",
X"c0",
X"80",
X"fc",
X"80",
X"c0",
X"00",
X"00",
X"00",
X"20",
X"60",
X"00",
X"f0",
X"fc",
X"fe",
X"66",
X"60",
X"30",
X"18",
X"0f",
X"1f",
X"3f",
X"3f",
X"7f",
X"7f",
X"3f",
X"1f",
X"00",
X"16",
X"2f",
X"2f",
X"20",
X"fc",
X"7c",
X"00",
X"00",
X"e0",
X"e0",
X"f0",
X"fe",
X"fc",
X"fc",
X"f8",
X"c0",
X"60",
X"20",
X"30",
X"3f",
X"3f",
X"3f",
X"3f",
X"3f",
X"3f",
X"3f",
X"1f",
X"2f",
X"2f",
X"2f",
X"0f",
X"07",
X"03",
X"00",
X"00",
X"f0",
X"90",
X"00",
X"08",
X"0c",
X"1c",
X"fc",
X"f8",
X"10",
X"f0",
X"f0",
X"f0",
X"f0",
X"e0",
X"c0",
X"e0",
X"0f",
X"0f",
X"07",
X"07",
X"07",
X"0f",
X"0f",
X"03",
X"01",
X"03",
X"01",
X"04",
X"07",
X"0f",
X"0f",
X"03",
X"f8",
X"f0",
X"e0",
X"f0",
X"b0",
X"80",
X"e0",
X"e0",
X"f8",
X"f0",
X"e0",
X"70",
X"b0",
X"80",
X"e0",
X"e0",
X"03",
X"3f",
X"7f",
X"19",
X"09",
X"09",
X"28",
X"5c",
X"00",
X"30",
X"70",
X"7f",
X"ff",
X"ff",
X"f7",
X"f3",
X"f8",
X"e0",
X"e0",
X"fc",
X"26",
X"30",
X"80",
X"10",
X"00",
X"18",
X"10",
X"00",
X"f8",
X"f8",
X"fe",
X"ff",
X"3e",
X"1e",
X"3f",
X"38",
X"30",
X"30",
X"00",
X"3a",
X"e7",
X"0f",
X"0f",
X"1f",
X"1f",
X"1f",
X"0f",
X"07",
X"78",
X"1e",
X"80",
X"fe",
X"7e",
X"7e",
X"7f",
X"7f",
X"ff",
X"fe",
X"fc",
X"c6",
X"8e",
X"ee",
X"ff",
X"ff",
X"3c",
X"3f",
X"1f",
X"0f",
X"07",
X"3f",
X"21",
X"20",
X"03",
X"00",
X"00",
X"0e",
X"07",
X"3f",
X"3f",
X"3f",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"fe",
X"fc",
X"70",
X"ff",
X"7f",
X"3f",
X"0e",
X"c0",
X"c0",
X"e0",
X"e0",
X"0f",
X"9f",
X"cf",
X"ff",
X"7f",
X"3f",
X"1e",
X"0e",
X"00",
X"80",
X"c8",
X"fe",
X"7f",
X"3f",
X"1e",
X"0e",
X"20",
X"c0",
X"80",
X"80",
X"00",
X"00",
X"00",
X"00",
X"e0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"03",
X"0f",
X"1f",
X"1f",
X"1c",
X"24",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"3f",
X"00",
X"04",
X"e6",
X"e0",
X"ff",
X"ff",
X"8f",
X"83",
X"0e",
X"1f",
X"1f",
X"1f",
X"1f",
X"03",
X"ff",
X"ff",
X"26",
X"26",
X"60",
X"78",
X"18",
X"0f",
X"7f",
X"ff",
X"3f",
X"3f",
X"7f",
X"7f",
X"1f",
X"00",
X"7e",
X"ff",
X"01",
X"21",
X"fe",
X"7a",
X"06",
X"fe",
X"fc",
X"fc",
X"ff",
X"ff",
X"fe",
X"fe",
X"fe",
X"de",
X"5c",
X"6c",
X"ff",
X"cf",
X"87",
X"07",
X"07",
X"0f",
X"1f",
X"1f",
X"ff",
X"ff",
X"fe",
X"fc",
X"f8",
X"b0",
X"60",
X"00",
X"f8",
X"f8",
X"f0",
X"b8",
X"f8",
X"f9",
X"fb",
X"ff",
X"28",
X"30",
X"18",
X"40",
X"00",
X"01",
X"03",
X"0f",
X"1f",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"c0",
X"80",
X"10",
X"ec",
X"e3",
X"e0",
X"e0",
X"e0",
X"c0",
X"80",
X"ff",
X"ff",
X"ff",
X"3f",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"13",
X"33",
X"30",
X"18",
X"04",
X"0f",
X"1f",
X"1f",
X"1f",
X"3f",
X"3f",
X"1f",
X"07",
X"09",
X"13",
X"17",
X"00",
X"10",
X"7e",
X"30",
X"e0",
X"f0",
X"f0",
X"e0",
X"ff",
X"ff",
X"fe",
X"ff",
X"fe",
X"fc",
X"f8",
X"e0",
X"1f",
X"1f",
X"0f",
X"0f",
X"0f",
X"1f",
X"1f",
X"1f",
X"17",
X"17",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"f0",
X"f8",
X"f8",
X"b8",
X"f8",
X"f8",
X"f8",
X"d0",
X"90",
X"18",
X"08",
X"40",
X"00",
X"00",
X"00",
X"3f",
X"ff",
X"ff",
X"ff",
X"f6",
X"c6",
X"84",
X"00",
X"30",
X"f0",
X"f0",
X"f1",
X"f6",
X"c6",
X"84",
X"00",
X"f0",
X"e0",
X"80",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"1f",
X"3f",
X"3f",
X"1f",
X"0f",
X"0f",
X"1f",
X"1f",
X"1f",
X"3f",
X"3e",
X"7c",
X"78",
X"f0",
X"e0",
X"f0",
X"f0",
X"f8",
X"f8",
X"b8",
X"f8",
X"f8",
X"f0",
X"b0",
X"90",
X"18",
X"08",
X"40",
X"00",
X"00",
X"00",
X"e0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f8",
X"f0",
X"c0",
X"e0",
X"fc",
X"fe",
X"ff",
X"7f",
X"03",
X"00",
X"1f",
X"1f",
X"1f",
X"3f",
X"3e",
X"3c",
X"38",
X"18",
X"00",
X"00",
X"10",
X"38",
X"3e",
X"3c",
X"38",
X"18",
X"00",
X"03",
X"07",
X"07",
X"0a",
X"0b",
X"0c",
X"00",
X"00",
X"00",
X"00",
X"07",
X"0f",
X"0f",
X"0f",
X"03",
X"00",
X"e0",
X"fc",
X"20",
X"20",
X"10",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"fc",
X"fe",
X"fc",
X"f8",
X"07",
X"07",
X"07",
X"1f",
X"1f",
X"3e",
X"21",
X"01",
X"07",
X"0f",
X"1b",
X"18",
X"10",
X"30",
X"21",
X"01",
X"e0",
X"e0",
X"e0",
X"f0",
X"f0",
X"e0",
X"c0",
X"e0",
X"a8",
X"fc",
X"f8",
X"00",
X"00",
X"00",
X"c0",
X"e0",
X"07",
X"0f",
X"0e",
X"14",
X"16",
X"18",
X"00",
X"3f",
X"00",
X"00",
X"0f",
X"1f",
X"1f",
X"1f",
X"07",
X"3c",
X"c0",
X"f8",
X"40",
X"40",
X"20",
X"78",
X"00",
X"c0",
X"00",
X"00",
X"e0",
X"f8",
X"fc",
X"f8",
X"f0",
X"c0",
X"3f",
X"0e",
X"0f",
X"1f",
X"3f",
X"7c",
X"70",
X"38",
X"fc",
X"ed",
X"c0",
X"00",
X"00",
X"60",
X"70",
X"38",
X"f0",
X"f8",
X"e4",
X"fc",
X"fc",
X"7c",
X"00",
X"00",
X"7e",
X"1e",
X"04",
X"0c",
X"0c",
X"0c",
X"00",
X"00",
X"07",
X"0f",
X"0e",
X"14",
X"16",
X"18",
X"00",
X"0f",
X"00",
X"00",
X"0f",
X"1f",
X"1f",
X"1f",
X"07",
X"0d",
X"1f",
X"1f",
X"1f",
X"1c",
X"0c",
X"07",
X"07",
X"07",
X"1e",
X"1c",
X"1e",
X"0f",
X"07",
X"00",
X"07",
X"07",
X"e0",
X"60",
X"f0",
X"70",
X"e0",
X"e0",
X"f0",
X"80",
X"60",
X"90",
X"00",
X"80",
X"00",
X"e0",
X"f0",
X"80",
X"07",
X"1f",
X"3f",
X"12",
X"13",
X"08",
X"1f",
X"31",
X"00",
X"10",
X"3f",
X"7f",
X"7f",
X"3f",
X"03",
X"0f",
X"c0",
X"f0",
X"40",
X"00",
X"30",
X"18",
X"c0",
X"f8",
X"00",
X"00",
X"e0",
X"f8",
X"fc",
X"f8",
X"b0",
X"38",
X"31",
X"39",
X"1f",
X"1f",
X"0f",
X"5f",
X"7e",
X"3c",
X"1f",
X"07",
X"00",
X"0e",
X"0f",
X"53",
X"7c",
X"3c",
X"f8",
X"f8",
X"f0",
X"e0",
X"e0",
X"c0",
X"00",
X"00",
X"f8",
X"f8",
X"f0",
X"00",
X"00",
X"80",
X"00",
X"00",
X"00",
X"e0",
X"fc",
X"27",
X"27",
X"11",
X"3e",
X"04",
X"07",
X"07",
X"03",
X"f7",
X"ff",
X"ff",
X"fe",
X"fc",
X"3f",
X"7f",
X"3f",
X"0f",
X"1f",
X"3f",
X"7f",
X"4f",
X"3e",
X"7f",
X"ff",
X"e2",
X"50",
X"38",
X"70",
X"40",
X"f8",
X"f9",
X"f9",
X"b7",
X"ff",
X"ff",
X"e0",
X"00",
X"e8",
X"71",
X"01",
X"4b",
X"03",
X"03",
X"00",
X"00",
X"07",
X"07",
X"0f",
X"3f",
X"3f",
X"3f",
X"26",
X"04",
X"05",
X"03",
X"01",
X"30",
X"30",
X"30",
X"26",
X"04",
X"f0",
X"f0",
X"f0",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"fe",
X"fc",
X"e0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"07",
X"07",
X"0f",
X"1f",
X"3f",
X"0f",
X"1c",
X"18",
X"05",
X"03",
X"01",
X"10",
X"30",
X"0c",
X"1c",
X"18",
X"e0",
X"e0",
X"e0",
X"e0",
X"c0",
X"80",
X"00",
X"00",
X"c0",
X"e0",
X"f0",
X"78",
X"18",
X"08",
X"00",
X"00",
X"07",
X"0f",
X"1f",
X"0f",
X"3f",
X"0f",
X"1c",
X"18",
X"07",
X"0f",
X"3e",
X"7c",
X"30",
X"0c",
X"1c",
X"18",
X"e0",
X"e0",
X"e0",
X"40",
X"c0",
X"80",
X"00",
X"00",
X"60",
X"60",
X"60",
X"80",
X"00",
X"00",
X"00",
X"00",
X"7f",
X"ff",
X"ff",
X"fb",
X"0f",
X"0f",
X"0f",
X"1f",
X"73",
X"f3",
X"f0",
X"f4",
X"f0",
X"f0",
X"70",
X"60",
X"3f",
X"7e",
X"7c",
X"7c",
X"3c",
X"3c",
X"fc",
X"fc",
X"00",
X"00",
X"00",
X"00",
X"3c",
X"3c",
X"fc",
X"fc",
X"60",
X"70",
X"18",
X"08",
X"0f",
X"1f",
X"3f",
X"7f",
X"7f",
X"7f",
X"1f",
X"07",
X"0b",
X"1b",
X"3b",
X"7b",
X"fc",
X"7c",
X"00",
X"20",
X"f0",
X"f8",
X"fc",
X"fe",
X"fc",
X"fc",
X"f8",
X"e0",
X"d0",
X"d8",
X"dc",
X"de",
X"0b",
X"0f",
X"1f",
X"1e",
X"3c",
X"3c",
X"3c",
X"7c",
X"c4",
X"e0",
X"e0",
X"40",
X"00",
X"3c",
X"3c",
X"7c",
X"1f",
X"3f",
X"0d",
X"07",
X"0f",
X"0e",
X"1c",
X"3c",
X"1d",
X"3c",
X"3a",
X"38",
X"30",
X"00",
X"1c",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"22",
X"55",
X"55",
X"55",
X"55",
X"55",
X"77",
X"22",
X"00",
X"07",
X"1f",
X"ff",
X"07",
X"1f",
X"0f",
X"06",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fb",
X"76",
X"00",
X"00",
X"cf",
X"07",
X"7f",
X"00",
X"00",
X"00",
X"20",
X"f8",
X"ff",
X"c3",
X"fd",
X"fe",
X"f0",
X"40",
X"00",
X"00",
X"3c",
X"fc",
X"fe",
X"e0",
X"00",
X"00",
X"40",
X"e0",
X"40",
X"40",
X"41",
X"41",
X"4f",
X"47",
X"40",
X"e0",
X"40",
X"3f",
X"3e",
X"3e",
X"30",
X"38",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"f8",
X"f8",
X"f8",
X"18",
X"38",
X"43",
X"46",
X"44",
X"40",
X"40",
X"40",
X"40",
X"40",
X"3c",
X"39",
X"3b",
X"3f",
X"00",
X"00",
X"00",
X"00",
X"80",
X"c0",
X"40",
X"00",
X"00",
X"00",
X"00",
X"00",
X"78",
X"38",
X"b8",
X"f8",
X"00",
X"00",
X"00",
X"00",
X"31",
X"30",
X"38",
X"7c",
X"7f",
X"ff",
X"ff",
X"fb",
X"3f",
X"3f",
X"0f",
X"77",
X"77",
X"f7",
X"f7",
X"f7",
X"10",
X"7e",
X"3e",
X"00",
X"1e",
X"fe",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"fe",
X"fa",
X"fa",
X"f3",
X"e7",
X"ff",
X"ff",
X"e3",
X"c3",
X"87",
X"48",
X"3c",
X"fc",
X"f0",
X"f8",
X"fc",
X"7c",
X"78",
X"38",
X"3c",
X"fc",
X"00",
X"ff",
X"c3",
X"83",
X"83",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"c3",
X"81",
X"81",
X"c3",
X"ff",
X"00",
X"1f",
X"1f",
X"0f",
X"07",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f0",
X"fb",
X"ff",
X"ff",
X"fe",
X"3e",
X"0c",
X"04",
X"00",
X"0b",
X"1f",
X"1f",
X"1e",
X"3e",
X"0c",
X"04",
X"1f",
X"1f",
X"0f",
X"0f",
X"07",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fb",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"03",
X"0f",
X"0f",
X"0f",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"18",
X"3c",
X"7e",
X"6e",
X"df",
X"df",
X"df",
X"00",
X"18",
X"3c",
X"7e",
X"76",
X"fb",
X"fb",
X"fb",
X"00",
X"18",
X"18",
X"3c",
X"3c",
X"3c",
X"3c",
X"1c",
X"00",
X"10",
X"10",
X"20",
X"20",
X"20",
X"20",
X"20",
X"00",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"00",
X"00",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"00",
X"08",
X"08",
X"04",
X"04",
X"04",
X"04",
X"04",
X"00",
X"10",
X"10",
X"38",
X"38",
X"38",
X"38",
X"38",
X"3c",
X"7e",
X"77",
X"fb",
X"9f",
X"5f",
X"8e",
X"20",
X"00",
X"18",
X"3c",
X"0e",
X"0e",
X"04",
X"00",
X"00",
X"5c",
X"2e",
X"8f",
X"3f",
X"7b",
X"77",
X"7e",
X"3c",
X"00",
X"00",
X"04",
X"06",
X"1e",
X"3c",
X"18",
X"00",
X"13",
X"4f",
X"3f",
X"bf",
X"3f",
X"7a",
X"f8",
X"f8",
X"00",
X"00",
X"01",
X"0a",
X"17",
X"0f",
X"2f",
X"1f",
X"00",
X"08",
X"05",
X"0f",
X"2f",
X"1d",
X"1c",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"05",
X"07",
X"0f",
X"07",
X"00",
X"00",
X"00",
X"00",
X"02",
X"0b",
X"07",
X"0f",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"08",
X"04",
X"04",
X"00",
X"60",
X"f0",
X"f8",
X"7c",
X"3e",
X"7e",
X"7f",
X"02",
X"02",
X"02",
X"05",
X"71",
X"7f",
X"7f",
X"7f",
X"3f",
X"5f",
X"7f",
X"3e",
X"0e",
X"0a",
X"51",
X"20",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"04",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0e",
X"1f",
X"02",
X"02",
X"00",
X"01",
X"13",
X"3f",
X"7f",
X"7f",
X"3f",
X"7f",
X"7f",
X"fe",
X"ec",
X"ca",
X"51",
X"20",
X"00",
X"40",
X"60",
X"70",
X"73",
X"27",
X"0f",
X"1f",
X"00",
X"40",
X"63",
X"77",
X"7c",
X"38",
X"f8",
X"e4",
X"00",
X"00",
X"00",
X"00",
X"03",
X"07",
X"0f",
X"1f",
X"00",
X"00",
X"03",
X"07",
X"0c",
X"18",
X"f8",
X"e4",
X"7f",
X"7f",
X"3f",
X"3f",
X"1f",
X"1f",
X"0f",
X"07",
X"03",
X"44",
X"28",
X"10",
X"08",
X"04",
X"03",
X"04",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"77",
X"77",
X"f5",
X"03",
X"07",
X"0f",
X"1f",
X"27",
X"7b",
X"78",
X"fb",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"ee",
X"ee",
X"af",
X"c0",
X"e0",
X"f0",
X"f8",
X"e4",
X"de",
X"1e",
X"df",
X"f1",
X"ff",
X"78",
X"00",
X"00",
X"18",
X"1c",
X"0e",
X"ff",
X"ff",
X"7f",
X"0f",
X"0f",
X"07",
X"03",
X"00",
X"8f",
X"ff",
X"1e",
X"00",
X"0c",
X"3e",
X"7e",
X"7c",
X"ff",
X"ff",
X"fe",
X"f0",
X"f0",
X"c0",
X"80",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"24",
X"24",
X"18",
X"00",
X"00",
X"00",
X"02",
X"41",
X"41",
X"61",
X"33",
X"06",
X"3c",
X"3c",
X"7e",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"3c",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"7f",
X"ff",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"63",
X"41",
X"c1",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"fe",
X"ff",
X"c0",
X"80",
X"00",
X"00",
X"8c",
X"fe",
X"fe",
X"f3",
X"ff",
X"ff",
X"ff",
X"78",
X"00",
X"00",
X"00",
X"00",
X"c1",
X"e3",
X"ff",
X"47",
X"0f",
X"0f",
X"0f",
X"07",
X"ff",
X"ff",
X"ff",
X"1e",
X"00",
X"20",
X"20",
X"40",
X"f1",
X"f9",
X"ff",
X"e2",
X"f0",
X"f0",
X"f0",
X"e0",
X"16",
X"1f",
X"3f",
X"7f",
X"3d",
X"1d",
X"3f",
X"1f",
X"16",
X"1f",
X"00",
X"00",
X"05",
X"0d",
X"3f",
X"1f",
X"80",
X"80",
X"c0",
X"e0",
X"f0",
X"f0",
X"f0",
X"f8",
X"80",
X"80",
X"00",
X"00",
X"00",
X"a0",
X"a0",
X"e0",
X"3c",
X"fa",
X"b1",
X"72",
X"f2",
X"db",
X"df",
X"5f",
X"00",
X"04",
X"4e",
X"8c",
X"0c",
X"7f",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"01",
X"01",
X"01",
X"06",
X"1e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"7f",
X"3f",
X"1f",
X"0f",
X"07",
X"03",
X"01",
X"00",
X"7c",
X"d6",
X"92",
X"ba",
X"ee",
X"fe",
X"38",
X"ff",
X"83",
X"29",
X"6d",
X"45",
X"11",
X"01",
X"c7",
X"00",
X"15",
X"3f",
X"62",
X"5f",
X"ff",
X"9f",
X"7d",
X"08",
X"08",
X"02",
X"1f",
X"22",
X"02",
X"02",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"08",
X"2f",
X"1e",
X"2f",
X"2f",
X"2f",
X"15",
X"0d",
X"0e",
X"10",
X"1e",
X"10",
X"50",
X"10",
X"08",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"1c",
X"3e",
X"7f",
X"ff",
X"ff",
X"fe",
X"7c",
X"38",
X"1c",
X"2a",
X"77",
X"ee",
X"dd",
X"aa",
X"74",
X"28",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"00",
X"ef",
X"ef",
X"ef",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"fe",
X"00",
X"ef",
X"ef",
X"ef",
X"00",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"7f",
X"5f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"68",
X"4e",
X"e0",
X"e0",
X"e0",
X"f0",
X"f8",
X"fc",
X"b8",
X"9e",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"7c",
X"3f",
X"5c",
X"39",
X"3b",
X"bb",
X"f9",
X"fc",
X"fe",
X"00",
X"23",
X"57",
X"4f",
X"57",
X"27",
X"c3",
X"21",
X"c0",
X"f0",
X"f0",
X"f0",
X"f0",
X"e0",
X"c0",
X"00",
X"00",
X"30",
X"70",
X"70",
X"f0",
X"e0",
X"c0",
X"00",
X"fe",
X"fc",
X"61",
X"0f",
X"ff",
X"fe",
X"f0",
X"e0",
X"13",
X"0f",
X"1e",
X"f0",
X"fc",
X"f8",
X"f0",
X"e0",
X"6e",
X"40",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"c0",
X"be",
X"90",
X"80",
X"c0",
X"c0",
X"80",
X"00",
X"00",
X"01",
X"01",
X"03",
X"03",
X"07",
X"7f",
X"7f",
X"3f",
X"01",
X"01",
X"03",
X"03",
X"07",
X"7f",
X"7d",
X"3d",
X"06",
X"07",
X"3f",
X"3c",
X"19",
X"7b",
X"7f",
X"3f",
X"06",
X"04",
X"30",
X"23",
X"06",
X"64",
X"60",
X"00",
X"3f",
X"7f",
X"7f",
X"1f",
X"3f",
X"3f",
X"07",
X"06",
X"00",
X"60",
X"60",
X"00",
X"20",
X"30",
X"04",
X"06",
X"03",
X"07",
X"0f",
X"0f",
X"0f",
X"0f",
X"07",
X"03",
X"00",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f8",
X"f8",
X"f8",
X"a0",
X"e1",
X"ff",
X"ff",
X"ff",
X"fe",
X"ff",
X"ff",
X"40",
X"01",
X"03",
X"03",
X"03",
X"0f",
X"0f",
X"0f",
X"1f",
X"1f",
X"1f",
X"0f",
X"07",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"e0",
X"f8",
X"f8",
X"f8",
X"ff",
X"fe",
X"f0",
X"c0",
X"e0",
X"fe",
X"ff",
X"7f",
X"03",
X"02",
X"00",
X"00",
X"01",
X"0f",
X"0f",
X"1f",
X"39",
X"33",
X"37",
X"7f",
X"01",
X"0d",
X"08",
X"00",
X"36",
X"2c",
X"08",
X"60",
X"7f",
X"3f",
X"3f",
X"3f",
X"1f",
X"0f",
X"0f",
X"01",
X"60",
X"00",
X"20",
X"30",
X"00",
X"08",
X"0d",
X"01",
X"00",
X"00",
X"03",
X"03",
X"47",
X"67",
X"77",
X"77",
X"01",
X"01",
X"03",
X"43",
X"67",
X"77",
X"7b",
X"78",
X"00",
X"00",
X"00",
X"00",
X"88",
X"98",
X"f8",
X"f0",
X"00",
X"00",
X"80",
X"84",
X"cc",
X"dc",
X"bc",
X"3c",
X"7e",
X"7f",
X"ff",
X"1f",
X"07",
X"30",
X"1c",
X"0c",
X"33",
X"07",
X"07",
X"e3",
X"38",
X"3f",
X"1c",
X"0c",
X"7e",
X"38",
X"f6",
X"ed",
X"df",
X"38",
X"70",
X"60",
X"98",
X"c7",
X"c8",
X"92",
X"30",
X"f8",
X"70",
X"60",
X"00",
X"00",
X"00",
X"03",
X"03",
X"47",
X"67",
X"77",
X"00",
X"01",
X"01",
X"03",
X"43",
X"67",
X"77",
X"7b",
X"00",
X"00",
X"00",
X"00",
X"00",
X"88",
X"98",
X"f8",
X"00",
X"00",
X"00",
X"80",
X"84",
X"cc",
X"dc",
X"bc",
X"77",
X"7e",
X"7f",
X"ff",
X"1f",
X"07",
X"70",
X"f0",
X"78",
X"33",
X"07",
X"07",
X"e3",
X"38",
X"7f",
X"f0",
X"f0",
X"7e",
X"38",
X"f6",
X"ed",
X"df",
X"38",
X"3c",
X"3c",
X"98",
X"c7",
X"c8",
X"92",
X"30",
X"f8",
X"3c",
X"03",
X"07",
X"0a",
X"1a",
X"1c",
X"1e",
X"0b",
X"08",
X"00",
X"10",
X"7f",
X"7f",
X"7f",
X"1f",
X"0f",
X"0f",
X"1c",
X"3f",
X"3f",
X"3d",
X"3f",
X"1f",
X"00",
X"00",
X"03",
X"33",
X"39",
X"3a",
X"38",
X"18",
X"00",
X"00",
X"00",
X"00",
X"04",
X"4c",
X"4e",
X"4e",
X"46",
X"6f",
X"10",
X"38",
X"3c",
X"74",
X"76",
X"76",
X"7e",
X"7d",
X"00",
X"1f",
X"3f",
X"3f",
X"4f",
X"5f",
X"7f",
X"7f",
X"00",
X"00",
X"11",
X"0a",
X"34",
X"2a",
X"51",
X"20",
X"7f",
X"67",
X"a3",
X"b0",
X"d8",
X"de",
X"dc",
X"c8",
X"7f",
X"67",
X"63",
X"70",
X"38",
X"3e",
X"7c",
X"b8",
X"7f",
X"7f",
X"7f",
X"1f",
X"47",
X"70",
X"70",
X"39",
X"51",
X"0a",
X"04",
X"ea",
X"79",
X"7f",
X"70",
X"39",
X"e8",
X"e8",
X"e0",
X"c0",
X"10",
X"70",
X"e0",
X"c0",
X"58",
X"38",
X"10",
X"30",
X"f0",
X"f0",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"20",
X"66",
X"66",
X"66",
X"62",
X"00",
X"08",
X"1c",
X"3c",
X"7a",
X"7a",
X"7a",
X"7e",
X"00",
X"00",
X"1f",
X"3f",
X"7f",
X"4f",
X"5f",
X"7f",
X"00",
X"00",
X"00",
X"11",
X"0a",
X"34",
X"2a",
X"51",
X"77",
X"7f",
X"3f",
X"b7",
X"b3",
X"db",
X"da",
X"d8",
X"7f",
X"7d",
X"3f",
X"37",
X"33",
X"3b",
X"3a",
X"78",
X"7f",
X"7f",
X"7f",
X"7f",
X"1f",
X"07",
X"70",
X"f0",
X"20",
X"51",
X"0a",
X"04",
X"ea",
X"39",
X"7f",
X"f0",
X"cc",
X"e8",
X"e8",
X"e0",
X"c0",
X"18",
X"7c",
X"3e",
X"bc",
X"58",
X"38",
X"10",
X"30",
X"f8",
X"fc",
X"3e",
X"03",
X"0f",
X"1f",
X"3f",
X"3b",
X"3f",
X"7f",
X"7f",
X"00",
X"00",
X"00",
X"06",
X"0e",
X"0c",
X"00",
X"00",
X"80",
X"f0",
X"f8",
X"fc",
X"fe",
X"fe",
X"ff",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"18",
X"7f",
X"7f",
X"7f",
X"7f",
X"ff",
X"0f",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f8",
X"3e",
X"3b",
X"18",
X"fe",
X"fb",
X"ff",
X"ff",
X"f6",
X"e0",
X"c0",
X"00",
X"10",
X"14",
X"10",
X"10",
X"38",
X"78",
X"f8",
X"30",
X"00",
X"03",
X"0f",
X"1f",
X"3f",
X"3b",
X"3f",
X"7f",
X"00",
X"00",
X"00",
X"00",
X"06",
X"0e",
X"0c",
X"00",
X"00",
X"c0",
X"f0",
X"f8",
X"fc",
X"fe",
X"fe",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"ff",
X"0f",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f8",
X"7e",
X"f3",
X"fe",
X"fe",
X"fb",
X"ff",
X"ff",
X"f6",
X"e0",
X"c0",
X"18",
X"10",
X"14",
X"10",
X"10",
X"38",
X"7c",
X"de",
X"00",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"08",
X"00",
X"0d",
X"1e",
X"1e",
X"1e",
X"1f",
X"0f",
X"07",
X"78",
X"f0",
X"f8",
X"e4",
X"c0",
X"ca",
X"ca",
X"c0",
X"78",
X"f0",
X"00",
X"1a",
X"3f",
X"35",
X"35",
X"3f",
X"0f",
X"1f",
X"9f",
X"ff",
X"ff",
X"7f",
X"74",
X"20",
X"00",
X"00",
X"80",
X"e0",
X"e0",
X"70",
X"73",
X"21",
X"e4",
X"ff",
X"fe",
X"fc",
X"9c",
X"1e",
X"00",
X"00",
X"1a",
X"07",
X"0c",
X"18",
X"78",
X"fe",
X"fc",
X"f0",
X"00",
X"01",
X"03",
X"03",
X"07",
X"03",
X"01",
X"00",
X"00",
X"01",
X"02",
X"00",
X"38",
X"7c",
X"7e",
X"3f",
X"00",
X"5f",
X"7f",
X"7f",
X"3f",
X"3f",
X"14",
X"00",
X"3f",
X"40",
X"60",
X"60",
X"20",
X"30",
X"13",
X"01",
X"c0",
X"e0",
X"f0",
X"30",
X"38",
X"3c",
X"3c",
X"fc",
X"c0",
X"e0",
X"30",
X"d0",
X"d0",
X"d0",
X"d0",
X"00",
X"07",
X"0f",
X"1f",
X"22",
X"20",
X"25",
X"25",
X"1f",
X"07",
X"0f",
X"02",
X"1d",
X"1f",
X"1a",
X"1a",
X"02",
X"fe",
X"fe",
X"7e",
X"3a",
X"02",
X"01",
X"41",
X"41",
X"38",
X"7c",
X"fc",
X"fc",
X"fc",
X"fe",
X"be",
X"be",
X"1f",
X"3f",
X"7e",
X"5c",
X"40",
X"80",
X"82",
X"82",
X"1c",
X"3e",
X"3f",
X"3f",
X"3f",
X"7f",
X"7d",
X"7d",
X"82",
X"80",
X"a0",
X"44",
X"43",
X"40",
X"21",
X"1e",
X"7d",
X"7f",
X"5f",
X"3b",
X"3c",
X"3f",
X"1e",
X"00",
X"1c",
X"3f",
X"3e",
X"3c",
X"40",
X"80",
X"82",
X"82",
X"1c",
X"3e",
X"3f",
X"1f",
X"3f",
X"7f",
X"7d",
X"7d",
X"00",
X"00",
X"80",
X"80",
X"92",
X"9d",
X"c7",
X"ef",
X"00",
X"00",
X"00",
X"60",
X"62",
X"65",
X"3f",
X"1f",
X"00",
X"23",
X"33",
X"3f",
X"3f",
X"7f",
X"7f",
X"7f",
X"70",
X"3c",
X"3c",
X"18",
X"00",
X"00",
X"02",
X"07",
X"fe",
X"f8",
X"a0",
X"00",
X"00",
X"00",
X"80",
X"80",
X"cf",
X"7a",
X"5a",
X"10",
X"00",
X"00",
X"c0",
X"80",
X"7e",
X"7f",
X"7d",
X"3f",
X"1e",
X"8f",
X"8f",
X"19",
X"85",
X"84",
X"86",
X"c6",
X"e7",
X"73",
X"73",
X"e1",
X"e0",
X"0e",
X"73",
X"f3",
X"f9",
X"f9",
X"f8",
X"70",
X"80",
X"4e",
X"77",
X"f3",
X"fb",
X"f9",
X"fa",
X"78",
X"0e",
X"66",
X"e2",
X"f6",
X"ff",
X"ff",
X"1f",
X"98",
X"11",
X"39",
X"7d",
X"39",
X"00",
X"00",
X"e0",
X"e7",
X"00",
X"00",
X"00",
X"04",
X"0f",
X"0f",
X"1f",
X"07",
X"00",
X"00",
X"07",
X"07",
X"16",
X"10",
X"00",
X"38",
X"f3",
X"e7",
X"ee",
X"ec",
X"cd",
X"cf",
X"cf",
X"df",
X"cf",
X"1f",
X"17",
X"10",
X"33",
X"30",
X"30",
X"20",
X"27",
X"3f",
X"3f",
X"78",
X"3c",
X"1f",
X"1f",
X"73",
X"38",
X"30",
X"40",
X"c7",
X"07",
X"66",
X"e0",
X"6c",
X"9f",
X"3e",
X"7c",
X"fc",
X"f8",
X"f8",
X"c0",
X"40",
X"60",
X"c0",
X"80",
X"04",
X"9e",
X"ff",
X"f0",
X"f8",
X"7f",
X"7e",
X"78",
X"01",
X"07",
X"1f",
X"3c",
X"7c",
X"24",
X"01",
X"07",
X"fe",
X"ff",
X"7f",
X"3f",
X"7f",
X"fc",
X"f8",
X"a0",
X"fe",
X"fc",
X"f0",
X"80",
X"00",
X"cf",
X"7a",
X"0a",
X"fe",
X"fc",
X"00",
X"00",
X"00",
X"7e",
X"7f",
X"7f",
X"3f",
X"1f",
X"8f",
X"8f",
X"18",
X"85",
X"86",
X"83",
X"c3",
X"e1",
X"70",
X"70",
X"e0",
X"9f",
X"3e",
X"7c",
X"f8",
X"f8",
X"3c",
X"18",
X"f8",
X"60",
X"c0",
X"80",
X"00",
X"98",
X"fc",
X"fe",
X"ff",
X"7f",
X"7f",
X"78",
X"01",
X"07",
X"13",
X"f1",
X"03",
X"24",
X"00",
X"07",
X"fe",
X"ff",
X"7f",
X"ff",
X"03",
X"00",
X"00",
X"1c",
X"1d",
X"1b",
X"c3",
X"e3",
X"e1",
X"03",
X"0f",
X"23",
X"62",
X"64",
X"3c",
X"1c",
X"1e",
X"e0",
X"cd",
X"1d",
X"4f",
X"ee",
X"ff",
X"3f",
X"3f",
X"1f",
X"3d",
X"6d",
X"4f",
X"ee",
X"f3",
X"20",
X"03",
X"3f",
X"3f",
X"00",
X"00",
X"70",
X"b8",
X"fc",
X"fc",
X"07",
X"07",
X"1f",
X"3f",
X"0f",
X"47",
X"03",
X"00",
X"07",
X"0f",
X"1f",
X"3f",
X"3e",
X"7c",
X"78",
X"78",
X"00",
X"00",
X"03",
X"07",
X"0f",
X"0f",
X"1f",
X"1f",
X"3f",
X"5c",
X"39",
X"3b",
X"bf",
X"ff",
X"fe",
X"fe",
X"00",
X"23",
X"57",
X"4f",
X"57",
X"2f",
X"df",
X"21",
X"c0",
X"c0",
X"80",
X"80",
X"80",
X"80",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"80",
X"80",
X"00",
X"00",
X"fe",
X"fc",
X"61",
X"0f",
X"7f",
X"3f",
X"1f",
X"1e",
X"23",
X"0f",
X"1e",
X"f0",
X"1c",
X"3f",
X"1f",
X"1e",
X"f0",
X"78",
X"e4",
X"c8",
X"cc",
X"be",
X"be",
X"3e",
X"00",
X"80",
X"18",
X"30",
X"34",
X"fe",
X"fe",
X"fe",
X"00",
X"01",
X"00",
X"07",
X"07",
X"07",
X"07",
X"1f",
X"00",
X"00",
X"01",
X"04",
X"06",
X"06",
X"07",
X"07",
X"00",
X"00",
X"0f",
X"3f",
X"3f",
X"0f",
X"00",
X"00",
X"0f",
X"3f",
X"7f",
X"f8",
X"f8",
X"7f",
X"3f",
X"0f",
X"78",
X"7c",
X"7e",
X"7f",
X"3f",
X"3f",
X"1b",
X"09",
X"1f",
X"1f",
X"1f",
X"0b",
X"01",
X"01",
X"00",
X"00",
X"0c",
X"00",
X"00",
X"00",
X"07",
X"7f",
X"7c",
X"00",
X"03",
X"1f",
X"3f",
X"3f",
X"78",
X"00",
X"03",
X"ff",
X"01",
X"e1",
X"71",
X"79",
X"3d",
X"3d",
X"1f",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"3f",
X"1f",
X"1b",
X"36",
X"30",
X"7f",
X"3f",
X"23",
X"27",
X"1f",
X"07",
X"0f",
X"1f",
X"7f",
X"3f",
X"f8",
X"f8",
X"f8",
X"b8",
X"18",
X"d8",
X"d8",
X"b8",
X"e0",
X"80",
X"80",
X"40",
X"e0",
X"e0",
X"e0",
X"c0",
X"01",
X"02",
X"04",
X"04",
X"08",
X"08",
X"10",
X"10",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"1f",
X"00",
X"0f",
X"13",
X"0d",
X"0d",
X"13",
X"0c",
X"20",
X"1f",
X"10",
X"0c",
X"12",
X"12",
X"2c",
X"3f",
X"3f",
X"00",
X"24",
X"00",
X"24",
X"00",
X"04",
X"00",
X"00",
X"37",
X"36",
X"36",
X"36",
X"16",
X"16",
X"12",
X"02",
X"0f",
X"41",
X"00",
X"88",
X"00",
X"44",
X"00",
X"00",
X"10",
X"7e",
X"ff",
X"ff",
X"f6",
X"76",
X"3a",
X"1a",
X"38",
X"7c",
X"fe",
X"fe",
X"3b",
X"03",
X"03",
X"03",
X"00",
X"00",
X"38",
X"04",
X"00",
X"00",
X"00",
X"00",
X"03",
X"33",
X"7b",
X"7f",
X"ff",
X"fb",
X"03",
X"03",
X"00",
X"00",
X"00",
X"38",
X"40",
X"00",
X"00",
X"00",
X"dc",
X"c0",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"c0",
X"fc",
X"a0",
X"80",
X"80",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"5f",
X"3f",
X"3f",
X"bb",
X"f8",
X"fe",
X"fe",
X"07",
X"27",
X"57",
X"4f",
X"57",
X"27",
X"c1",
X"21",
X"1f",
X"0f",
X"0f",
X"1f",
X"1f",
X"1e",
X"38",
X"30",
X"1d",
X"0f",
X"0f",
X"1f",
X"1f",
X"1e",
X"38",
X"30",
X"00",
X"20",
X"60",
X"60",
X"70",
X"f0",
X"f8",
X"f8",
X"00",
X"00",
X"38",
X"10",
X"4c",
X"18",
X"86",
X"24",
X"f8",
X"fc",
X"fc",
X"7e",
X"7e",
X"3e",
X"1f",
X"07",
X"00",
X"42",
X"0a",
X"40",
X"10",
X"02",
X"08",
X"02",
X"00",
X"c0",
X"70",
X"b8",
X"f4",
X"f2",
X"f5",
X"7b",
X"00",
X"00",
X"80",
X"40",
X"08",
X"0c",
X"0a",
X"84",
X"00",
X"df",
X"10",
X"ff",
X"df",
X"ff",
X"ff",
X"f9",
X"00",
X"00",
X"cf",
X"20",
X"20",
X"20",
X"26",
X"2e",
X"1f",
X"1f",
X"3e",
X"fc",
X"f8",
X"f0",
X"c0",
X"00",
X"e0",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f8",
X"fc",
X"fe",
X"ff",
X"ff",
X"df",
X"df",
X"00",
X"2f",
X"23",
X"21",
X"20",
X"20",
X"00",
X"00",
X"00",
X"c1",
X"f1",
X"79",
X"7d",
X"3d",
X"3f",
X"1f",
X"03",
X"c1",
X"b1",
X"59",
X"6d",
X"35",
X"3b",
X"1f",
X"03",
X"02",
X"06",
X"0e",
X"0e",
X"1e",
X"1e",
X"3e",
X"3e",
X"00",
X"02",
X"00",
X"08",
X"02",
X"00",
X"28",
X"00",
X"3e",
X"3e",
X"3e",
X"3e",
X"1e",
X"1e",
X"0e",
X"02",
X"04",
X"10",
X"02",
X"10",
X"04",
X"00",
X"0a",
X"00",
X"c1",
X"f1",
X"79",
X"7d",
X"3d",
X"3f",
X"1f",
X"03",
X"c1",
X"b1",
X"59",
X"6d",
X"35",
X"3b",
X"1f",
X"03",
X"7c",
X"00",
X"00",
X"ff",
X"c3",
X"7f",
X"1f",
X"03",
X"00",
X"0f",
X"1f",
X"ff",
X"fc",
X"63",
X"1f",
X"03",
X"ff",
X"ff",
X"7c",
X"00",
X"00",
X"7c",
X"ff",
X"ff",
X"00",
X"00",
X"fe",
X"c6",
X"c6",
X"fe",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"04",
X"0c",
X"18",
X"30",
X"00",
X"00",
X"00",
X"06",
X"06",
X"0c",
X"18",
X"70",
X"60",
X"ff",
X"ff",
X"00",
X"04",
X"04",
X"04",
X"08",
X"08",
X"00",
X"00",
X"06",
X"06",
X"04",
X"04",
X"08",
X"08",
X"08",
X"10",
X"10",
X"00",
X"00",
X"10",
X"10",
X"08",
X"08",
X"10",
X"30",
X"30",
X"30",
X"30",
X"10",
X"08",
X"7f",
X"3f",
X"3f",
X"3e",
X"1f",
X"0f",
X"03",
X"00",
X"00",
X"00",
X"01",
X"03",
X"01",
X"00",
X"00",
X"00",
X"03",
X"0f",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"03",
X"0e",
X"f8",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"22",
X"65",
X"25",
X"25",
X"25",
X"25",
X"77",
X"72",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"62",
X"95",
X"15",
X"25",
X"45",
X"85",
X"f7",
X"f2",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"a2",
X"a5",
X"a5",
X"a5",
X"f5",
X"f5",
X"27",
X"22",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f2",
X"85",
X"85",
X"e5",
X"15",
X"15",
X"f7",
X"e2",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"62",
X"95",
X"55",
X"65",
X"b5",
X"95",
X"97",
X"62",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"20",
X"50",
X"50",
X"50",
X"50",
X"50",
X"70",
X"20",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"e6",
X"66",
X"66",
X"66",
X"67",
X"f3",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"5e",
X"59",
X"59",
X"59",
X"5e",
X"d8",
X"98",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"38",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"04",
X"08",
X"00",
X"38",
X"4c",
X"c6",
X"c6",
X"c6",
X"64",
X"38",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"38",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"c6",
X"0e",
X"3c",
X"78",
X"e0",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7e",
X"0c",
X"18",
X"3c",
X"06",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1c",
X"3c",
X"6c",
X"cc",
X"fe",
X"0c",
X"0c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fc",
X"c0",
X"fc",
X"06",
X"06",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"3c",
X"60",
X"c0",
X"fc",
X"c6",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fe",
X"c6",
X"0c",
X"18",
X"30",
X"30",
X"30",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"c6",
X"c6",
X"7c",
X"c6",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"c6",
X"c6",
X"7e",
X"06",
X"0c",
X"78",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"38",
X"6c",
X"c6",
X"c6",
X"fe",
X"c6",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fc",
X"c6",
X"c6",
X"fc",
X"c6",
X"c6",
X"fc",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"3c",
X"66",
X"c0",
X"c0",
X"c0",
X"66",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"f8",
X"cc",
X"c6",
X"c6",
X"c6",
X"cc",
X"f8",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fe",
X"c0",
X"c0",
X"fc",
X"c0",
X"c0",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fe",
X"c0",
X"c0",
X"fc",
X"c0",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"3e",
X"60",
X"c0",
X"ce",
X"c6",
X"66",
X"3e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"c6",
X"c6",
X"fe",
X"c6",
X"c6",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1e",
X"06",
X"06",
X"06",
X"c6",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"cc",
X"d8",
X"f0",
X"f8",
X"dc",
X"ce",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"60",
X"60",
X"60",
X"60",
X"60",
X"60",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"ee",
X"fe",
X"fe",
X"d6",
X"c6",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"e6",
X"f6",
X"fe",
X"de",
X"ce",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"c6",
X"c6",
X"c6",
X"c6",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fc",
X"c6",
X"c6",
X"c6",
X"fc",
X"c0",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7c",
X"c6",
X"c6",
X"c6",
X"de",
X"cc",
X"7a",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fc",
X"c6",
X"c6",
X"ce",
X"f8",
X"dc",
X"ce",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"78",
X"cc",
X"c0",
X"7c",
X"06",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7e",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"c6",
X"c6",
X"c6",
X"c6",
X"c6",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"c6",
X"c6",
X"ee",
X"7c",
X"38",
X"10",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"c6",
X"d6",
X"fe",
X"fe",
X"ee",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"c6",
X"ee",
X"7c",
X"38",
X"7c",
X"ee",
X"c6",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"66",
X"66",
X"66",
X"3c",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fe",
X"0e",
X"1c",
X"38",
X"70",
X"e0",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"7e",
X"7e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"44",
X"28",
X"10",
X"28",
X"44",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"18",
X"3c",
X"3c",
X"3c",
X"18",
X"18",
X"00",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"ff",
X"e3",
X"c1",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"00",
X"1c",
X"3e",
X"80",
X"80",
X"80",
X"c1",
X"e3",
X"ff",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"3e",
X"1c",
X"00",
X"00",
X"ff",
X"38",
X"7c",
X"7c",
X"7c",
X"7c",
X"7c",
X"38",
X"00",
X"08",
X"04",
X"04",
X"04",
X"04",
X"04",
X"08",
X"00",
X"03",
X"06",
X"0c",
X"0c",
X"08",
X"08",
X"04",
X"03",
X"03",
X"05",
X"0b",
X"0b",
X"0f",
X"0f",
X"07",
X"03",
X"01",
X"02",
X"04",
X"08",
X"10",
X"20",
X"40",
X"80",
X"01",
X"03",
X"07",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"07",
X"38",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"07",
X"3f",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"e0",
X"1c",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"e0",
X"fc",
X"ff",
X"80",
X"40",
X"20",
X"10",
X"08",
X"04",
X"02",
X"01",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"ff",
X"04",
X"0e",
X"0e",
X"0e",
X"6e",
X"64",
X"60",
X"60",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"07",
X"0f",
X"1f",
X"1f",
X"7f",
X"ff",
X"ff",
X"7f",
X"07",
X"08",
X"10",
X"00",
X"60",
X"80",
X"80",
X"40",
X"03",
X"07",
X"1f",
X"3f",
X"3f",
X"3f",
X"79",
X"f7",
X"03",
X"04",
X"18",
X"20",
X"20",
X"20",
X"46",
X"88",
X"c0",
X"e0",
X"f0",
X"f4",
X"fe",
X"bf",
X"df",
X"ff",
X"c0",
X"20",
X"10",
X"14",
X"0a",
X"41",
X"21",
X"01",
X"90",
X"b8",
X"f8",
X"fa",
X"ff",
X"ff",
X"ff",
X"fe",
X"90",
X"a8",
X"48",
X"0a",
X"05",
X"01",
X"01",
X"02",
X"3b",
X"1d",
X"0e",
X"0f",
X"07",
X"00",
X"00",
X"00",
X"24",
X"12",
X"09",
X"08",
X"07",
X"00",
X"00",
X"00",
X"ff",
X"bf",
X"1c",
X"c0",
X"f3",
X"ff",
X"7e",
X"1c",
X"00",
X"40",
X"e3",
X"3f",
X"0c",
X"81",
X"62",
X"1c",
X"bf",
X"7f",
X"3d",
X"83",
X"c7",
X"ff",
X"ff",
X"3c",
X"40",
X"80",
X"c2",
X"7c",
X"38",
X"00",
X"c3",
X"3c",
X"fc",
X"fe",
X"ff",
X"fe",
X"fe",
X"f8",
X"60",
X"00",
X"04",
X"02",
X"01",
X"00",
X"06",
X"98",
X"60",
X"00",
X"c0",
X"20",
X"10",
X"10",
X"10",
X"10",
X"20",
X"c0",
X"c0",
X"e0",
X"f0",
X"f0",
X"f0",
X"f0",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"3f",
X"7f",
X"e0",
X"c0",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1c",
X"3e",
X"88",
X"9c",
X"88",
X"80",
X"80",
X"80",
X"80",
X"80",
X"7f",
X"7f",
X"7f",
X"3e",
X"1c",
X"00",
X"00",
X"00",
X"fe",
X"fe",
X"fe",
X"fe",
X"fe",
X"fe",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"08",
X"14",
X"24",
X"c4",
X"03",
X"40",
X"a1",
X"26",
X"00",
X"08",
X"18",
X"38",
X"fc",
X"bf",
X"5e",
X"d9",
X"ff",
X"ff",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"7f",
X"80",
X"80",
X"98",
X"9c",
X"8c",
X"80",
X"80",
X"00",
X"7f",
X"7f",
X"67",
X"67",
X"7f",
X"7f",
X"7f",
X"ff",
X"01",
X"01",
X"ff",
X"10",
X"10",
X"10",
X"ff",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"01",
X"01",
X"01",
X"ff",
X"10",
X"10",
X"10",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"01",
X"01",
X"19",
X"1d",
X"0d",
X"01",
X"01",
X"00",
X"ff",
X"ff",
X"e7",
X"e7",
X"ff",
X"ff",
X"ff",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"3f",
X"7f",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"3f",
X"60",
X"40",
X"c0",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"3c",
X"80",
X"80",
X"80",
X"80",
X"80",
X"81",
X"42",
X"3c",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"82",
X"7c",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"7c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"83",
X"ff",
X"f8",
X"fc",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"f8",
X"04",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"3c",
X"01",
X"01",
X"01",
X"01",
X"01",
X"81",
X"42",
X"3c",
X"00",
X"08",
X"08",
X"08",
X"10",
X"10",
X"10",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"7f",
X"7f",
X"78",
X"73",
X"73",
X"73",
X"7f",
X"7f",
X"80",
X"a0",
X"87",
X"8f",
X"8e",
X"8e",
X"86",
X"00",
X"ff",
X"ff",
X"3f",
X"9f",
X"9f",
X"9f",
X"1f",
X"fe",
X"01",
X"05",
X"c1",
X"e1",
X"71",
X"71",
X"f1",
X"7e",
X"7e",
X"7f",
X"7e",
X"7e",
X"7f",
X"7f",
X"ff",
X"81",
X"81",
X"80",
X"81",
X"81",
X"a0",
X"80",
X"ff",
X"7f",
X"7f",
X"ff",
X"7f",
X"7f",
X"ff",
X"ff",
X"ff",
X"f1",
X"c1",
X"c1",
X"81",
X"c1",
X"c5",
X"01",
X"ff",
X"7f",
X"80",
X"a0",
X"80",
X"80",
X"80",
X"80",
X"80",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"01",
X"05",
X"01",
X"01",
X"01",
X"01",
X"01",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"80",
X"a0",
X"80",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7f",
X"01",
X"01",
X"01",
X"01",
X"01",
X"05",
X"01",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"00",
X"00",
X"00",
X"00",
X"fc",
X"fe",
X"07",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"38",
X"7c",
X"11",
X"39",
X"11",
X"01",
X"01",
X"01",
X"01",
X"01",
X"fe",
X"fe",
X"fe",
X"7c",
X"38",
X"00",
X"00",
X"00",
X"ef",
X"28",
X"28",
X"28",
X"28",
X"28",
X"ef",
X"00",
X"20",
X"e7",
X"e7",
X"e7",
X"e7",
X"e7",
X"ef",
X"00",
X"fe",
X"82",
X"82",
X"82",
X"82",
X"82",
X"fe",
X"00",
X"02",
X"7e",
X"7e",
X"7e",
X"7e",
X"7e",
X"fe",
X"00",
X"80",
X"80",
X"80",
X"98",
X"9c",
X"8c",
X"80",
X"7f",
X"7f",
X"7f",
X"7f",
X"67",
X"67",
X"7f",
X"7f",
X"7f",
X"ff",
X"ff",
X"83",
X"f3",
X"f3",
X"f3",
X"f3",
X"f3",
X"ff",
X"80",
X"fc",
X"8c",
X"8c",
X"8c",
X"8c",
X"8c",
X"ff",
X"ff",
X"f0",
X"f6",
X"f6",
X"f6",
X"f6",
X"f6",
X"ff",
X"00",
X"0f",
X"09",
X"09",
X"09",
X"09",
X"09",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"01",
X"57",
X"2f",
X"57",
X"2f",
X"57",
X"ff",
X"01",
X"ff",
X"a9",
X"d1",
X"a9",
X"d1",
X"a9",
X"f3",
X"f3",
X"f3",
X"f3",
X"f3",
X"f3",
X"ff",
X"3f",
X"8c",
X"8c",
X"8c",
X"8c",
X"8c",
X"8c",
X"ff",
X"3f",
X"f6",
X"f6",
X"f6",
X"f6",
X"f6",
X"f6",
X"ff",
X"ff",
X"09",
X"09",
X"09",
X"09",
X"09",
X"09",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"2f",
X"57",
X"2f",
X"57",
X"2f",
X"57",
X"ff",
X"fc",
X"d1",
X"a9",
X"d1",
X"a9",
X"d1",
X"a9",
X"ff",
X"fc",
X"3c",
X"3c",
X"3c",
X"3c",
X"3c",
X"3c",
X"3c",
X"3c",
X"23",
X"23",
X"23",
X"23",
X"23",
X"23",
X"23",
X"23",
X"fb",
X"fb",
X"fb",
X"fb",
X"fb",
X"fb",
X"fb",
X"fb",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"04",
X"bc",
X"5c",
X"bc",
X"5c",
X"bc",
X"5c",
X"bc",
X"5c",
X"44",
X"a4",
X"44",
X"a4",
X"44",
X"a4",
X"44",
X"a4",
X"1f",
X"20",
X"40",
X"40",
X"80",
X"80",
X"80",
X"81",
X"1f",
X"3f",
X"7f",
X"7f",
X"ff",
X"ff",
X"ff",
X"fe",
X"ff",
X"80",
X"80",
X"c0",
X"ff",
X"ff",
X"fe",
X"fe",
X"ff",
X"7f",
X"7f",
X"3f",
X"00",
X"00",
X"01",
X"01",
X"ff",
X"7f",
X"7f",
X"ff",
X"ff",
X"07",
X"03",
X"03",
X"ff",
X"80",
X"80",
X"00",
X"00",
X"f8",
X"fc",
X"fc",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"81",
X"c3",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"3c",
X"00",
X"f8",
X"fc",
X"fe",
X"fe",
X"e3",
X"c1",
X"81",
X"81",
X"f8",
X"04",
X"02",
X"02",
X"1d",
X"3f",
X"7f",
X"7f",
X"83",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7f",
X"1f",
X"fc",
X"80",
X"80",
X"80",
X"80",
X"80",
X"60",
X"1f",
X"fc",
X"fc",
X"fc",
X"fc",
X"fe",
X"fe",
X"ff",
X"ff",
X"03",
X"03",
X"03",
X"03",
X"01",
X"01",
X"00",
X"ff",
X"01",
X"01",
X"01",
X"01",
X"03",
X"03",
X"07",
X"ff",
X"fe",
X"fe",
X"fe",
X"fe",
X"fc",
X"fc",
X"f8",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"81",
X"c1",
X"e3",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"7f",
X"3f",
X"1d",
X"01",
X"01",
X"01",
X"03",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fb",
X"b5",
X"ce",
X"80",
X"80",
X"80",
X"80",
X"80",
X"84",
X"ca",
X"b1",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"df",
X"ad",
X"73",
X"01",
X"01",
X"01",
X"01",
X"01",
X"21",
X"53",
X"8d",
X"77",
X"77",
X"77",
X"77",
X"77",
X"77",
X"77",
X"77",
X"00",
X"00",
X"00",
X"00",
X"77",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"77",
X"77",
X"77",
X"77",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"77",
X"77",
X"77",
X"77",
X"77",
X"01",
X"01",
X"01",
X"19",
X"1d",
X"0d",
X"01",
X"fe",
X"ff",
X"ff",
X"ff",
X"e7",
X"e7",
X"ff",
X"ff",
X"fe",
X"20",
X"78",
X"7f",
X"fe",
X"fe",
X"fe",
X"fe",
X"fe",
X"00",
X"21",
X"21",
X"41",
X"41",
X"41",
X"41",
X"41",
X"04",
X"9a",
X"fa",
X"fd",
X"fd",
X"fd",
X"fd",
X"fd",
X"00",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"7e",
X"38",
X"21",
X"00",
X"01",
X"00",
X"01",
X"00",
X"21",
X"21",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"fa",
X"8a",
X"84",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"02",
X"04",
X"00",
X"10",
X"00",
X"40",
X"80",
X"00",
X"01",
X"01",
X"06",
X"08",
X"18",
X"20",
X"20",
X"c0",
X"0b",
X"0b",
X"3b",
X"0b",
X"fb",
X"0b",
X"0b",
X"0a",
X"04",
X"04",
X"c4",
X"f4",
X"f4",
X"04",
X"04",
X"05",
X"90",
X"10",
X"1f",
X"10",
X"1f",
X"10",
X"10",
X"90",
X"70",
X"f0",
X"f0",
X"ff",
X"ff",
X"f0",
X"f0",
X"70",
X"3f",
X"78",
X"e7",
X"cf",
X"58",
X"58",
X"50",
X"90",
X"c0",
X"87",
X"18",
X"b0",
X"e7",
X"e7",
X"ef",
X"ef",
X"b0",
X"fc",
X"e2",
X"c1",
X"c1",
X"83",
X"8f",
X"7e",
X"6f",
X"43",
X"5d",
X"3f",
X"3f",
X"7f",
X"7f",
X"ff",
X"fe",
X"03",
X"0f",
X"91",
X"70",
X"60",
X"20",
X"31",
X"03",
X"ff",
X"f1",
X"6e",
X"cf",
X"df",
X"ff",
X"ff",
X"3f",
X"3f",
X"1d",
X"39",
X"7b",
X"f3",
X"86",
X"fe",
X"fd",
X"fb",
X"fb",
X"f7",
X"f7",
X"0f",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"ff",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"80",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"03",
X"03",
X"ff",
X"fe",
X"03",
X"03",
X"03",
X"03",
X"ff",
X"ff",
X"03",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"3c",
X"fc",
X"fc",
X"fc",
X"fc",
X"fc",
X"04",
X"04",
X"23",
X"f3",
X"0b",
X"0b",
X"0b",
X"07",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"ff",
X"ff",
X"03",
X"ff",
X"ff",
X"ff",
X"03",
X"03",
X"03",
X"03",
X"ff",
X"03",
X"03",
X"03",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"00",
X"00",
X"fc",
X"fc",
X"fe",
X"fe",
X"fe",
X"02",
X"fe",
X"fe",
X"07",
X"07",
X"03",
X"03",
X"03",
X"ff",
X"03",
X"03",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"04",
X"04",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"aa",
X"d5",
X"aa",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"d5",
X"aa",
X"d5",
X"80",
X"80",
X"ff",
X"03",
X"03",
X"ab",
X"57",
X"ab",
X"ff",
X"ff",
X"fe",
X"ff",
X"ff",
X"57",
X"ab",
X"57",
X"03",
X"03",
X"fe",
X"00",
X"55",
X"aa",
X"55",
X"ff",
X"ff",
X"ff",
X"00",
X"ff",
X"aa",
X"55",
X"aa",
X"00",
X"00",
X"ff",
X"00",
X"04",
X"54",
X"ac",
X"5c",
X"fc",
X"fc",
X"fc",
X"3c",
X"ff",
X"af",
X"57",
X"ab",
X"0b",
X"0b",
X"f3",
X"23",
X"3f",
X"3f",
X"3f",
X"3f",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"7c",
X"7c",
X"78",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"1f",
X"0f",
X"0f",
X"07",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"fc",
X"fc",
X"f8",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"07",
X"1f",
X"3f",
X"ff",
X"7f",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"e1",
X"f9",
X"fd",
X"ff",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"f0",
X"10",
X"10",
X"10",
X"10",
X"10",
X"10",
X"ff",
X"00",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"1f",
X"10",
X"10",
X"10",
X"10",
X"10",
X"10",
X"ff",
X"00",
X"0f",
X"0f",
X"0f",
X"0f",
X"0f",
X"0f",
X"0f",
X"92",
X"92",
X"92",
X"fe",
X"fe",
X"00",
X"00",
X"00",
X"48",
X"48",
X"6c",
X"00",
X"00",
X"00",
X"fe",
X"00",
X"0a",
X"0a",
X"3a",
X"0a",
X"fb",
X"0b",
X"0b",
X"0b",
X"05",
X"05",
X"c5",
X"f5",
X"f4",
X"04",
X"04",
X"04",
X"90",
X"90",
X"9f",
X"90",
X"9f",
X"90",
X"90",
X"90",
X"70",
X"70",
X"70",
X"7f",
X"7f",
X"70",
X"70",
X"70",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"08",
X"88",
X"91",
X"d1",
X"53",
X"53",
X"73",
X"3f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"be",
X"ce",
X"00",
X"00",
X"07",
X"0f",
X"0c",
X"1b",
X"1b",
X"1b",
X"00",
X"00",
X"00",
X"00",
X"03",
X"04",
X"04",
X"04",
X"00",
X"00",
X"e0",
X"f0",
X"f0",
X"f8",
X"f8",
X"f8",
X"00",
X"00",
X"60",
X"30",
X"30",
X"98",
X"98",
X"98",
X"1b",
X"1b",
X"1b",
X"1b",
X"1b",
X"0f",
X"0f",
X"07",
X"04",
X"04",
X"04",
X"04",
X"04",
X"03",
X"00",
X"00",
X"f8",
X"f8",
X"f8",
X"f8",
X"f8",
X"f0",
X"f0",
X"e0",
X"98",
X"98",
X"98",
X"98",
X"98",
X"30",
X"30",
X"60",
X"f1",
X"11",
X"11",
X"1f",
X"10",
X"10",
X"10",
X"ff",
X"0f",
X"ef",
X"ef",
X"ef",
X"ef",
X"ef",
X"ef",
X"e0",
X"1f",
X"10",
X"10",
X"f0",
X"10",
X"10",
X"10",
X"ff",
X"e0",
X"ef",
X"ef",
X"ef",
X"ef",
X"ef",
X"ef",
X"0f",
X"7f",
X"bf",
X"df",
X"ef",
X"f0",
X"f0",
X"f0",
X"f0",
X"80",
X"40",
X"20",
X"10",
X"0f",
X"0f",
X"0f",
X"0f",
X"f0",
X"f0",
X"f0",
X"f0",
X"ff",
X"ff",
X"ff",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"1f",
X"3f",
X"7f",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"01",
X"03",
X"07",
X"0f",
X"ff",
X"ff",
X"ff",
X"ff",
X"0f",
X"0f",
X"0f",
X"0f",
X"f7",
X"fb",
X"fd",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"18",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"1f",
X"3f",
X"7f",
X"7f",
X"7f",
X"ff",
X"ff",
X"ff",
X"1f",
X"20",
X"40",
X"40",
X"40",
X"80",
X"82",
X"82",
X"ff",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"3f",
X"1e",
X"82",
X"80",
X"a0",
X"44",
X"43",
X"40",
X"21",
X"1e",
X"f8",
X"fc",
X"fe",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"f8",
X"04",
X"02",
X"02",
X"02",
X"01",
X"41",
X"41",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"fe",
X"fc",
X"78",
X"41",
X"01",
X"05",
X"22",
X"c2",
X"02",
X"84",
X"78",
X"7f",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"de",
X"61",
X"61",
X"61",
X"71",
X"5e",
X"7f",
X"61",
X"61",
X"df",
X"df",
X"df",
X"df",
X"ff",
X"c1",
X"df",
X"80",
X"80",
X"c0",
X"f0",
X"bf",
X"8f",
X"81",
X"7e",
X"7f",
X"7f",
X"ff",
X"3f",
X"4f",
X"71",
X"7f",
X"ff",
X"61",
X"61",
X"c1",
X"c1",
X"81",
X"81",
X"83",
X"fe",
X"df",
X"df",
X"bf",
X"bf",
X"7f",
X"7f",
X"7f",
X"7f",
X"00",
X"00",
X"03",
X"0f",
X"1f",
X"3f",
X"7f",
X"7f",
X"00",
X"00",
X"03",
X"0c",
X"10",
X"20",
X"40",
X"40",
X"00",
X"00",
X"c0",
X"f0",
X"f8",
X"fc",
X"fe",
X"fe",
X"00",
X"00",
X"c0",
X"30",
X"08",
X"04",
X"02",
X"02",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"7f",
X"7f",
X"7f",
X"3f",
X"3f",
X"1f",
X"0f",
X"07",
X"40",
X"40",
X"40",
X"20",
X"30",
X"1c",
X"0f",
X"07",
X"fe",
X"fe",
X"fe",
X"fc",
X"fc",
X"f8",
X"f0",
X"f0",
X"02",
X"02",
X"02",
X"04",
X"0c",
X"38",
X"f0",
X"f0",
X"0f",
X"0f",
X"0f",
X"0f",
X"0f",
X"0f",
X"07",
X"0f",
X"08",
X"08",
X"08",
X"08",
X"08",
X"0c",
X"05",
X"0a",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"f0",
X"e0",
X"f0",
X"10",
X"50",
X"50",
X"50",
X"50",
X"30",
X"a0",
X"50",
X"81",
X"c1",
X"a3",
X"a3",
X"9d",
X"81",
X"81",
X"81",
X"00",
X"41",
X"22",
X"22",
X"1c",
X"00",
X"00",
X"00",
X"e3",
X"f7",
X"c1",
X"c1",
X"c1",
X"c1",
X"f7",
X"e3",
X"e3",
X"14",
X"3e",
X"3e",
X"3e",
X"3e",
X"14",
X"e3",
X"00",
X"00",
X"07",
X"0f",
X"0c",
X"1b",
X"1b",
X"1b",
X"ff",
X"ff",
X"f8",
X"f0",
X"f0",
X"e0",
X"e0",
X"e0",
X"00",
X"00",
X"e0",
X"f0",
X"f0",
X"f8",
X"f8",
X"f8",
X"ff",
X"ff",
X"7f",
X"3f",
X"3f",
X"9f",
X"9f",
X"9f",
X"1b",
X"1b",
X"1b",
X"1b",
X"1b",
X"0f",
X"0f",
X"07",
X"e0",
X"e0",
X"e0",
X"e0",
X"e0",
X"f3",
X"f0",
X"f8",
X"f8",
X"f8",
X"f8",
X"f8",
X"f8",
X"f0",
X"f0",
X"e0",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"3f",
X"3f",
X"7f",
X"e0",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"70",
X"1f",
X"10",
X"70",
X"7f",
X"7f",
X"7f",
X"07",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"03",
X"f8",
X"00",
X"03",
X"fb",
X"fb",
X"fb",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"ff",
X"ef",
X"7c",
X"7b",
X"76",
X"75",
X"75",
X"77",
X"17",
X"67",
X"ff",
X"df",
X"ef",
X"af",
X"af",
X"6f",
X"ef",
X"e7",
X"3b",
X"fb",
X"7b",
X"fb",
X"fb",
X"f3",
X"f8",
X"f3",
X"1f",
X"1f",
X"3f",
X"3f",
X"70",
X"63",
X"e7",
X"e5",
X"0f",
X"0f",
X"1f",
X"1f",
X"3f",
X"3c",
X"78",
X"7a",
X"f0",
X"f0",
X"f8",
X"f8",
X"0c",
X"c4",
X"e4",
X"a6",
X"f8",
X"f8",
X"fc",
X"fc",
X"fe",
X"3e",
X"1e",
X"5f",
X"e9",
X"e9",
X"e9",
X"ef",
X"e2",
X"e3",
X"f0",
X"ff",
X"76",
X"76",
X"76",
X"70",
X"7d",
X"7c",
X"7f",
X"7f",
X"96",
X"96",
X"96",
X"f6",
X"46",
X"c6",
X"0e",
X"fe",
X"6f",
X"6f",
X"6f",
X"0f",
X"bf",
X"3f",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"7e",
X"3c",
X"3c",
X"7e",
X"7e",
X"ff",
X"ff",
X"ff",
X"42",
X"00",
X"3c",
X"42",
X"99",
X"a1",
X"a1",
X"99",
X"42",
X"3c",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0f",
X"1f",
X"1f",
X"3f",
X"3f",
X"7f",
X"7f",
X"7f",
X"f0",
X"e0",
X"e0",
X"c0",
X"c0",
X"80",
X"80",
X"80",
X"f0",
X"f8",
X"f8",
X"fc",
X"fc",
X"fe",
X"fe",
X"fe",
X"0f",
X"07",
X"07",
X"03",
X"03",
X"01",
X"01",
X"01",
X"7f",
X"7f",
X"3f",
X"3f",
X"3f",
X"3f",
X"1f",
X"1f",
X"80",
X"80",
X"c0",
X"c0",
X"e0",
X"f8",
X"fe",
X"ff",
X"fe",
X"ff",
X"ff",
X"ff",
X"fc",
X"fc",
X"fe",
X"fe",
X"ff",
X"7f",
X"1f",
X"07",
X"03",
X"03",
X"01",
X"81",
X"7f",
X"7f",
X"7f",
X"3f",
X"3f",
X"3f",
X"3f",
X"1f",
X"80",
X"80",
X"80",
X"c0",
X"c0",
X"e0",
X"e0",
X"f0",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"01",
X"01",
X"01",
X"03",
X"03",
X"07",
X"07",
X"0f",
X"1f",
X"0f",
X"0f",
X"07",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"fc",
X"fc",
X"f8",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"7e",
X"7e",
X"7e",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"01",
X"01",
X"01",
X"03",
X"03",
X"07",
X"07",
X"0f",
X"fe",
X"fe",
X"fe",
X"fe",
X"ff",
X"ff",
X"ff",
X"ff",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"ff",
X"ff",
X"ff",
X"ff",
X"fc",
X"fe",
X"fe",
X"7e",
X"ff",
X"03",
X"03",
X"03",
X"03",
X"03",
X"03",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"80",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"01",
X"01",
X"01",
X"03",
X"07",
X"03",
X"01",
X"01",
X"7e",
X"7e",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"3f",
X"3f",
X"3f",
X"3f",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"7e",
X"7c",
X"7c",
X"78",
X"00",
X"00",
X"00",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"fe",
X"fe",
X"ff",
X"ff",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"7f",
X"7f",
X"3f",
X"3f",
X"3f",
X"3f",
X"1f",
X"1f",
X"80",
X"80",
X"c0",
X"c0",
X"e0",
X"f8",
X"fe",
X"ff",
X"3f",
X"bf",
X"ff",
X"ff",
X"fc",
X"fc",
X"fe",
X"fe",
X"ff",
X"7f",
X"1f",
X"07",
X"03",
X"03",
X"01",
X"81",
X"7f",
X"7f",
X"7e",
X"7e",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"7e",
X"7e",
X"7e",
X"7e",
X"7f",
X"7f",
X"7f",
X"7f",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"81",
X"c3",
X"c3",
X"e7",
X"e7",
X"ff",
X"ff",
X"ff",
X"7e",
X"3c",
X"3c",
X"18",
X"18",
X"00",
X"00",
X"00",
X"0f",
X"43",
X"5b",
X"53",
X"31",
X"19",
X"0f",
X"07",
X"f2",
X"fe",
X"fe",
X"ff",
X"ff",
X"ef",
X"f7",
X"f8",
X"c1",
X"c3",
X"c6",
X"84",
X"fc",
X"fc",
X"0e",
X"02",
X"bf",
X"be",
X"bd",
X"7b",
X"7b",
X"07",
X"f3",
X"fd",
X"10",
X"20",
X"22",
X"ba",
X"e6",
X"e1",
X"c0",
X"c0",
X"ff",
X"ff",
X"ff",
X"67",
X"59",
X"9e",
X"bf",
X"bf",
X"20",
X"a6",
X"54",
X"26",
X"20",
X"c6",
X"54",
X"26",
X"20",
X"e6",
X"54",
X"26",
X"21",
X"06",
X"54",
X"26",
X"20",
X"85",
X"01",
X"44",
X"20",
X"86",
X"54",
X"48",
X"20",
X"9a",
X"01",
X"49",
X"20",
X"a5",
X"c9",
X"46",
X"20",
X"ba",
X"c9",
X"4a",
X"20",
X"a6",
X"0a",
X"d0",
X"d1",
X"d8",
X"d8",
X"de",
X"d1",
X"d0",
X"da",
X"de",
X"d1",
X"20",
X"c6",
X"0a",
X"d2",
X"d3",
X"db",
X"db",
X"db",
X"d9",
X"db",
X"dc",
X"db",
X"df",
X"20",
X"e6",
X"0a",
X"d4",
X"d5",
X"d4",
X"d9",
X"db",
X"e2",
X"d4",
X"da",
X"db",
X"e0",
X"21",
X"06",
X"0a",
X"d6",
X"d7",
X"d6",
X"d7",
X"e1",
X"26",
X"d6",
X"dd",
X"e1",
X"e1",
X"21",
X"26",
X"14",
X"d0",
X"e8",
X"d1",
X"d0",
X"d1",
X"de",
X"d1",
X"d8",
X"d0",
X"d1",
X"26",
X"de",
X"d1",
X"de",
X"d1",
X"d0",
X"d1",
X"d0",
X"d1",
X"26",
X"21",
X"46",
X"14",
X"db",
X"42",
X"42",
X"db",
X"42",
X"db",
X"42",
X"db",
X"db",
X"42",
X"26",
X"db",
X"42",
X"db",
X"42",
X"db",
X"42",
X"db",
X"42",
X"26",
X"21",
X"66",
X"46",
X"db",
X"21",
X"6c",
X"0e",
X"df",
X"db",
X"db",
X"db",
X"26",
X"db",
X"df",
X"db",
X"df",
X"db",
X"db",
X"e4",
X"e5",
X"26",
X"21",
X"86",
X"14",
X"db",
X"db",
X"db",
X"de",
X"43",
X"db",
X"e0",
X"db",
X"db",
X"db",
X"26",
X"db",
X"e3",
X"db",
X"e0",
X"db",
X"db",
X"e6",
X"e3",
X"26",
X"21",
X"a6",
X"14",
X"db",
X"db",
X"db",
X"db",
X"42",
X"db",
X"db",
X"db",
X"d4",
X"d9",
X"26",
X"db",
X"d9",
X"db",
X"db",
X"d4",
X"d9",
X"d4",
X"d9",
X"e7",
X"21",
X"c5",
X"16",
X"5f",
X"95",
X"95",
X"95",
X"95",
X"95",
X"95",
X"95",
X"95",
X"97",
X"98",
X"78",
X"95",
X"96",
X"95",
X"95",
X"97",
X"98",
X"97",
X"98",
X"95",
X"7a",
X"21",
X"ed",
X"0e",
X"cf",
X"01",
X"09",
X"08",
X"05",
X"24",
X"17",
X"12",
X"17",
X"1d",
X"0e",
X"17",
X"0d",
X"18",
X"22",
X"4b",
X"0d",
X"01",
X"24",
X"19",
X"15",
X"0a",
X"22",
X"0e",
X"1b",
X"24",
X"10",
X"0a",
X"16",
X"0e",
X"22",
X"8b",
X"0d",
X"02",
X"24",
X"19",
X"15",
X"0a",
X"22",
X"0e",
X"1b",
X"24",
X"10",
X"0a",
X"16",
X"0e",
X"22",
X"ec",
X"04",
X"1d",
X"18",
X"19",
X"28",
X"22",
X"f6",
X"01",
X"00",
X"23",
X"c9",
X"56",
X"55",
X"23",
X"e2",
X"04",
X"99",
X"aa",
X"aa",
X"aa",
X"23",
X"ea",
X"04",
X"99",
X"aa",
X"aa",
X"aa",
X"00",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff"
);
	
	begin
	
	process(clock)
	begin
		if(rising_edge(clock)) then
			q_a <= rom(address_a);
			q_b <= rom(address_b);
		end if;
	end process;

end rtl;
