library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is

	port
	(
		address		: in natural range 0 to 32767;
		clock		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
	
end entity;

architecture rtl of rom is

	-- Build a 2-D array type for the RoM
	-- subtype word_t is std_logic_vector(7 downto 0);
	-- type memory_t is array(32767 downto 0) of word_t;
	subtype word_t is std_logic_vector(0 to 7);
	type memory_t is array(0 to 32767) of word_t;
		
	-- function init_rom
	-- 	return memory_t is
	-- 	variable tmp : memory_t := (others => (others => '0'));
	-- 	begin
	-- 		for addr_pos in 0 to 32767 loop
	-- 			-- Initialize each address with the address itself
	-- 			tmp(addr_pos) := std_logic_vector(to_unsigned(addr_pos, 8));
	-- 		end loop;
	-- 	return tmp;
	-- end init_rom;
	
	-- Declare the ROM signal and specify a default value.	Quartus II
	-- will create a memory initialization file (.mif) based on the 
	-- default value.
	-- signal rom : memory_t := init_rom;
	signal rom : memory_t := 
(
X"78",
X"d8",
X"a9",
X"10",
X"8d",
X"00",
X"20",
X"a2",
X"ff",
X"9a",
X"ad",
X"02",
X"20",
X"10",
X"fb",
X"ad",
X"02",
X"20",
X"10",
X"fb",
X"a0",
X"fe",
X"a2",
X"05",
X"bd",
X"d7",
X"07",
X"c9",
X"0a",
X"b0",
X"0c",
X"ca",
X"10",
X"f6",
X"ad",
X"ff",
X"07",
X"c9",
X"a5",
X"d0",
X"02",
X"a0",
X"d6",
X"20",
X"cc",
X"90",
X"8d",
X"11",
X"40",
X"8d",
X"70",
X"07",
X"a9",
X"a5",
X"8d",
X"ff",
X"07",
X"8d",
X"a7",
X"07",
X"a9",
X"0f",
X"8d",
X"15",
X"40",
X"a9",
X"06",
X"8d",
X"01",
X"20",
X"20",
X"20",
X"82",
X"20",
X"19",
X"8e",
X"ee",
X"74",
X"07",
X"ad",
X"78",
X"07",
X"09",
X"80",
X"20",
X"ed",
X"8e",
X"4c",
X"57",
X"80",
X"01",
X"a4",
X"c8",
X"ec",
X"10",
X"00",
X"41",
X"41",
X"4c",
X"34",
X"3c",
X"44",
X"54",
X"68",
X"7c",
X"a8",
X"bf",
X"de",
X"ef",
X"03",
X"8c",
X"8c",
X"8c",
X"8d",
X"03",
X"03",
X"03",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"8d",
X"00",
X"40",
X"ad",
X"78",
X"07",
X"29",
X"7f",
X"8d",
X"78",
X"07",
X"29",
X"7e",
X"8d",
X"00",
X"20",
X"ad",
X"79",
X"07",
X"29",
X"e6",
X"ac",
X"74",
X"07",
X"d0",
X"05",
X"ad",
X"79",
X"07",
X"09",
X"1e",
X"8d",
X"79",
X"07",
X"29",
X"e7",
X"8d",
X"01",
X"20",
X"ae",
X"02",
X"20",
X"a9",
X"00",
X"20",
X"e6",
X"8e",
X"8d",
X"03",
X"20",
X"a9",
X"02",
X"8d",
X"14",
X"40",
X"ae",
X"73",
X"07",
X"bd",
X"5a",
X"80",
X"85",
X"00",
X"bd",
X"6d",
X"80",
X"85",
X"01",
X"20",
X"dd",
X"8e",
X"a0",
X"00",
X"ae",
X"73",
X"07",
X"e0",
X"06",
X"d0",
X"01",
X"c8",
X"be",
X"80",
X"80",
X"a9",
X"00",
X"9d",
X"00",
X"03",
X"9d",
X"01",
X"03",
X"8d",
X"73",
X"07",
X"ad",
X"79",
X"07",
X"8d",
X"01",
X"20",
X"20",
X"d0",
X"f2",
X"20",
X"5c",
X"8e",
X"20",
X"82",
X"81",
X"20",
X"97",
X"8f",
X"ad",
X"76",
X"07",
X"4a",
X"b0",
X"25",
X"ad",
X"47",
X"07",
X"f0",
X"05",
X"ce",
X"47",
X"07",
X"d0",
X"19",
X"a2",
X"14",
X"ce",
X"7f",
X"07",
X"10",
X"07",
X"a9",
X"14",
X"8d",
X"7f",
X"07",
X"a2",
X"23",
X"bd",
X"80",
X"07",
X"f0",
X"03",
X"de",
X"80",
X"07",
X"ca",
X"10",
X"f5",
X"e6",
X"09",
X"a2",
X"00",
X"a0",
X"07",
X"ad",
X"a7",
X"07",
X"29",
X"02",
X"85",
X"00",
X"ad",
X"a8",
X"07",
X"29",
X"02",
X"45",
X"00",
X"18",
X"f0",
X"01",
X"38",
X"7e",
X"a7",
X"07",
X"e8",
X"88",
X"d0",
X"f9",
X"ad",
X"22",
X"07",
X"f0",
X"1f",
X"ad",
X"02",
X"20",
X"29",
X"40",
X"d0",
X"f9",
X"ad",
X"76",
X"07",
X"4a",
X"b0",
X"06",
X"20",
X"23",
X"82",
X"20",
X"c6",
X"81",
X"ad",
X"02",
X"20",
X"29",
X"40",
X"f0",
X"f9",
X"a0",
X"14",
X"88",
X"d0",
X"fd",
X"ad",
X"3f",
X"07",
X"8d",
X"05",
X"20",
X"ad",
X"40",
X"07",
X"8d",
X"05",
X"20",
X"ad",
X"78",
X"07",
X"48",
X"8d",
X"00",
X"20",
X"ad",
X"76",
X"07",
X"4a",
X"b0",
X"03",
X"20",
X"12",
X"82",
X"ad",
X"02",
X"20",
X"68",
X"09",
X"80",
X"8d",
X"00",
X"20",
X"40",
X"ad",
X"70",
X"07",
X"c9",
X"02",
X"f0",
X"0b",
X"c9",
X"01",
X"d0",
X"38",
X"ad",
X"72",
X"07",
X"c9",
X"03",
X"d0",
X"31",
X"ad",
X"77",
X"07",
X"f0",
X"04",
X"ce",
X"77",
X"07",
X"60",
X"ad",
X"fc",
X"06",
X"29",
X"10",
X"f0",
X"19",
X"ad",
X"76",
X"07",
X"29",
X"80",
X"d0",
X"1a",
X"a9",
X"2b",
X"8d",
X"77",
X"07",
X"ad",
X"76",
X"07",
X"a8",
X"c8",
X"84",
X"fa",
X"49",
X"01",
X"09",
X"80",
X"d0",
X"05",
X"ad",
X"76",
X"07",
X"29",
X"7f",
X"8d",
X"76",
X"07",
X"60",
X"ac",
X"4e",
X"07",
X"a9",
X"28",
X"85",
X"00",
X"a2",
X"0e",
X"bd",
X"e4",
X"06",
X"c5",
X"00",
X"90",
X"0f",
X"ac",
X"e0",
X"06",
X"18",
X"79",
X"e1",
X"06",
X"90",
X"03",
X"18",
X"65",
X"00",
X"9d",
X"e4",
X"06",
X"ca",
X"10",
X"e7",
X"ae",
X"e0",
X"06",
X"e8",
X"e0",
X"03",
X"d0",
X"02",
X"a2",
X"00",
X"8e",
X"e0",
X"06",
X"a2",
X"08",
X"a0",
X"02",
X"b9",
X"e9",
X"06",
X"9d",
X"f1",
X"06",
X"18",
X"69",
X"08",
X"9d",
X"f2",
X"06",
X"18",
X"69",
X"08",
X"9d",
X"f3",
X"06",
X"ca",
X"ca",
X"ca",
X"88",
X"10",
X"e8",
X"60",
X"ad",
X"70",
X"07",
X"20",
X"04",
X"8e",
X"31",
X"82",
X"dc",
X"ae",
X"8b",
X"83",
X"18",
X"92",
X"a0",
X"00",
X"2c",
X"a0",
X"04",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"c8",
X"c8",
X"c8",
X"c8",
X"d0",
X"f7",
X"60",
X"ad",
X"72",
X"07",
X"20",
X"04",
X"8e",
X"cf",
X"8f",
X"67",
X"85",
X"61",
X"90",
X"45",
X"82",
X"04",
X"20",
X"73",
X"01",
X"00",
X"00",
X"a0",
X"00",
X"ad",
X"fc",
X"06",
X"0d",
X"fd",
X"06",
X"c9",
X"10",
X"f0",
X"04",
X"c9",
X"90",
X"d0",
X"03",
X"4c",
X"d8",
X"82",
X"c9",
X"20",
X"f0",
X"1a",
X"ae",
X"a2",
X"07",
X"d0",
X"0b",
X"8d",
X"80",
X"07",
X"20",
X"6b",
X"83",
X"b0",
X"60",
X"4c",
X"c0",
X"82",
X"ae",
X"fc",
X"07",
X"f0",
X"4a",
X"c9",
X"40",
X"d0",
X"46",
X"c8",
X"ad",
X"a2",
X"07",
X"f0",
X"4e",
X"a9",
X"18",
X"8d",
X"a2",
X"07",
X"ad",
X"80",
X"07",
X"d0",
X"36",
X"a9",
X"10",
X"8d",
X"80",
X"07",
X"c0",
X"01",
X"f0",
X"0e",
X"ad",
X"7a",
X"07",
X"49",
X"01",
X"8d",
X"7a",
X"07",
X"20",
X"25",
X"83",
X"4c",
X"bb",
X"82",
X"ae",
X"6b",
X"07",
X"e8",
X"8a",
X"29",
X"07",
X"8d",
X"6b",
X"07",
X"20",
X"0e",
X"83",
X"bd",
X"3f",
X"82",
X"9d",
X"00",
X"03",
X"e8",
X"e0",
X"06",
X"30",
X"f5",
X"ac",
X"5f",
X"07",
X"c8",
X"8c",
X"04",
X"03",
X"a9",
X"00",
X"8d",
X"fc",
X"06",
X"20",
X"ea",
X"ae",
X"a5",
X"0e",
X"c9",
X"06",
X"d0",
X"44",
X"a9",
X"00",
X"8d",
X"70",
X"07",
X"8d",
X"72",
X"07",
X"8d",
X"22",
X"07",
X"ee",
X"74",
X"07",
X"60",
X"ac",
X"a2",
X"07",
X"f0",
X"ec",
X"0a",
X"90",
X"06",
X"ad",
X"fd",
X"07",
X"20",
X"0e",
X"83",
X"20",
X"03",
X"9c",
X"ee",
X"5d",
X"07",
X"ee",
X"64",
X"07",
X"ee",
X"57",
X"07",
X"ee",
X"70",
X"07",
X"ad",
X"fc",
X"07",
X"8d",
X"6a",
X"07",
X"a9",
X"00",
X"8d",
X"72",
X"07",
X"8d",
X"a2",
X"07",
X"a2",
X"17",
X"a9",
X"00",
X"9d",
X"dd",
X"07",
X"ca",
X"10",
X"fa",
X"60",
X"8d",
X"5f",
X"07",
X"8d",
X"66",
X"07",
X"a2",
X"00",
X"8e",
X"60",
X"07",
X"8e",
X"67",
X"07",
X"60",
X"07",
X"22",
X"49",
X"83",
X"ce",
X"24",
X"24",
X"00",
X"a0",
X"07",
X"b9",
X"1d",
X"83",
X"99",
X"00",
X"03",
X"88",
X"10",
X"f7",
X"ad",
X"7a",
X"07",
X"f0",
X"0a",
X"a9",
X"24",
X"8d",
X"04",
X"03",
X"a9",
X"ce",
X"8d",
X"06",
X"03",
X"60",
X"01",
X"80",
X"02",
X"81",
X"41",
X"80",
X"01",
X"42",
X"c2",
X"02",
X"80",
X"41",
X"c1",
X"41",
X"c1",
X"01",
X"c1",
X"01",
X"02",
X"80",
X"00",
X"9b",
X"10",
X"18",
X"05",
X"2c",
X"20",
X"24",
X"15",
X"5a",
X"10",
X"20",
X"28",
X"30",
X"20",
X"10",
X"80",
X"20",
X"30",
X"30",
X"01",
X"ff",
X"00",
X"ae",
X"17",
X"07",
X"ad",
X"18",
X"07",
X"d0",
X"0d",
X"e8",
X"ee",
X"17",
X"07",
X"38",
X"bd",
X"54",
X"83",
X"8d",
X"18",
X"07",
X"f0",
X"0a",
X"bd",
X"3f",
X"83",
X"8d",
X"fc",
X"06",
X"ce",
X"18",
X"07",
X"18",
X"60",
X"20",
X"a0",
X"83",
X"ad",
X"72",
X"07",
X"f0",
X"07",
X"a2",
X"00",
X"86",
X"08",
X"20",
X"47",
X"c0",
X"20",
X"2a",
X"f1",
X"4c",
X"e9",
X"ee",
X"ad",
X"72",
X"07",
X"20",
X"04",
X"8e",
X"ec",
X"cf",
X"b0",
X"83",
X"bd",
X"83",
X"f6",
X"83",
X"61",
X"84",
X"ae",
X"1b",
X"07",
X"e8",
X"86",
X"34",
X"a9",
X"08",
X"85",
X"fc",
X"4c",
X"4e",
X"87",
X"a0",
X"00",
X"84",
X"35",
X"a5",
X"6d",
X"c5",
X"34",
X"d0",
X"06",
X"a5",
X"86",
X"c9",
X"60",
X"b0",
X"03",
X"e6",
X"35",
X"c8",
X"98",
X"20",
X"e6",
X"b0",
X"ad",
X"1a",
X"07",
X"c5",
X"34",
X"f0",
X"16",
X"ad",
X"68",
X"07",
X"18",
X"69",
X"80",
X"8d",
X"68",
X"07",
X"a9",
X"01",
X"69",
X"00",
X"a8",
X"20",
X"c4",
X"af",
X"20",
X"6f",
X"af",
X"e6",
X"35",
X"a5",
X"35",
X"f0",
X"68",
X"60",
X"ad",
X"49",
X"07",
X"d0",
X"48",
X"ad",
X"19",
X"07",
X"f0",
X"18",
X"c9",
X"09",
X"b0",
X"3f",
X"ac",
X"5f",
X"07",
X"c0",
X"07",
X"d0",
X"09",
X"c9",
X"03",
X"90",
X"34",
X"e9",
X"01",
X"4c",
X"18",
X"84",
X"c9",
X"02",
X"90",
X"2b",
X"a8",
X"d0",
X"08",
X"ad",
X"53",
X"07",
X"f0",
X"14",
X"c8",
X"d0",
X"11",
X"c8",
X"ad",
X"5f",
X"07",
X"c9",
X"07",
X"f0",
X"09",
X"88",
X"c0",
X"04",
X"b0",
X"26",
X"c0",
X"03",
X"b0",
X"0f",
X"c0",
X"03",
X"d0",
X"04",
X"a9",
X"04",
X"85",
X"fc",
X"98",
X"18",
X"69",
X"0c",
X"8d",
X"73",
X"07",
X"ad",
X"49",
X"07",
X"18",
X"69",
X"04",
X"8d",
X"49",
X"07",
X"ad",
X"19",
X"07",
X"69",
X"00",
X"8d",
X"19",
X"07",
X"c9",
X"07",
X"90",
X"08",
X"a9",
X"06",
X"8d",
X"a1",
X"07",
X"ee",
X"72",
X"07",
X"60",
X"ad",
X"a1",
X"07",
X"d0",
X"20",
X"ac",
X"5f",
X"07",
X"c0",
X"07",
X"b0",
X"1a",
X"a9",
X"00",
X"8d",
X"60",
X"07",
X"8d",
X"5c",
X"07",
X"8d",
X"72",
X"07",
X"ee",
X"5f",
X"07",
X"20",
X"03",
X"9c",
X"ee",
X"57",
X"07",
X"a9",
X"01",
X"8d",
X"70",
X"07",
X"60",
X"ad",
X"fc",
X"06",
X"0d",
X"fd",
X"06",
X"29",
X"40",
X"f0",
X"0d",
X"a9",
X"01",
X"8d",
X"fc",
X"07",
X"a9",
X"ff",
X"8d",
X"5a",
X"07",
X"20",
X"48",
X"92",
X"60",
X"ff",
X"ff",
X"f6",
X"fb",
X"f7",
X"fb",
X"f8",
X"fb",
X"f9",
X"fb",
X"fa",
X"fb",
X"f6",
X"50",
X"f7",
X"50",
X"f8",
X"50",
X"f9",
X"50",
X"fa",
X"50",
X"fd",
X"fe",
X"ff",
X"41",
X"42",
X"44",
X"45",
X"48",
X"31",
X"32",
X"34",
X"35",
X"38",
X"00",
X"bd",
X"10",
X"01",
X"f0",
X"be",
X"c9",
X"0b",
X"90",
X"05",
X"a9",
X"0b",
X"9d",
X"10",
X"01",
X"a8",
X"bd",
X"2c",
X"01",
X"d0",
X"04",
X"9d",
X"10",
X"01",
X"60",
X"de",
X"2c",
X"01",
X"c9",
X"2b",
X"d0",
X"1e",
X"c0",
X"0b",
X"d0",
X"07",
X"ee",
X"5a",
X"07",
X"a9",
X"40",
X"85",
X"fe",
X"b9",
X"b7",
X"84",
X"4a",
X"4a",
X"4a",
X"4a",
X"aa",
X"b9",
X"b7",
X"84",
X"29",
X"0f",
X"9d",
X"34",
X"01",
X"20",
X"27",
X"bc",
X"bc",
X"e5",
X"06",
X"b5",
X"16",
X"c9",
X"12",
X"f0",
X"22",
X"c9",
X"0d",
X"f0",
X"1e",
X"c9",
X"05",
X"f0",
X"12",
X"c9",
X"0a",
X"f0",
X"16",
X"c9",
X"0b",
X"f0",
X"12",
X"c9",
X"09",
X"b0",
X"06",
X"b5",
X"1e",
X"c9",
X"02",
X"b0",
X"08",
X"ae",
X"ee",
X"03",
X"bc",
X"ec",
X"06",
X"a6",
X"08",
X"bd",
X"1e",
X"01",
X"c9",
X"18",
X"90",
X"05",
X"e9",
X"01",
X"9d",
X"1e",
X"01",
X"bd",
X"1e",
X"01",
X"e9",
X"08",
X"20",
X"c1",
X"e5",
X"bd",
X"17",
X"01",
X"99",
X"03",
X"02",
X"18",
X"69",
X"08",
X"99",
X"07",
X"02",
X"a9",
X"02",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"bd",
X"10",
X"01",
X"0a",
X"aa",
X"bd",
X"9f",
X"84",
X"99",
X"01",
X"02",
X"bd",
X"a0",
X"84",
X"99",
X"05",
X"02",
X"a6",
X"08",
X"60",
X"ad",
X"3c",
X"07",
X"20",
X"04",
X"8e",
X"8b",
X"85",
X"9b",
X"85",
X"52",
X"86",
X"5a",
X"86",
X"93",
X"86",
X"9d",
X"88",
X"a8",
X"86",
X"9d",
X"88",
X"e6",
X"86",
X"bf",
X"85",
X"e3",
X"85",
X"43",
X"86",
X"ff",
X"86",
X"32",
X"87",
X"49",
X"87",
X"20",
X"20",
X"82",
X"20",
X"19",
X"8e",
X"ad",
X"70",
X"07",
X"f0",
X"32",
X"a2",
X"03",
X"4c",
X"c5",
X"85",
X"ad",
X"44",
X"07",
X"48",
X"ad",
X"56",
X"07",
X"48",
X"a9",
X"00",
X"8d",
X"56",
X"07",
X"a9",
X"02",
X"8d",
X"44",
X"07",
X"20",
X"f1",
X"85",
X"68",
X"8d",
X"56",
X"07",
X"68",
X"8d",
X"44",
X"07",
X"4c",
X"45",
X"87",
X"01",
X"02",
X"03",
X"04",
X"ac",
X"4e",
X"07",
X"be",
X"bb",
X"85",
X"8e",
X"73",
X"07",
X"4c",
X"45",
X"87",
X"00",
X"09",
X"0a",
X"04",
X"22",
X"22",
X"0f",
X"0f",
X"0f",
X"22",
X"0f",
X"0f",
X"22",
X"16",
X"27",
X"18",
X"22",
X"30",
X"27",
X"19",
X"22",
X"37",
X"27",
X"16",
X"ac",
X"44",
X"07",
X"f0",
X"06",
X"b9",
X"c7",
X"85",
X"8d",
X"73",
X"07",
X"ee",
X"3c",
X"07",
X"ae",
X"00",
X"03",
X"a0",
X"00",
X"ad",
X"53",
X"07",
X"f0",
X"02",
X"a0",
X"04",
X"ad",
X"56",
X"07",
X"c9",
X"02",
X"d0",
X"02",
X"a0",
X"08",
X"a9",
X"03",
X"85",
X"00",
X"b9",
X"d7",
X"85",
X"9d",
X"04",
X"03",
X"c8",
X"e8",
X"c6",
X"00",
X"10",
X"f4",
X"ae",
X"00",
X"03",
X"ac",
X"44",
X"07",
X"d0",
X"03",
X"ac",
X"4e",
X"07",
X"b9",
X"cf",
X"85",
X"9d",
X"04",
X"03",
X"a9",
X"3f",
X"9d",
X"01",
X"03",
X"a9",
X"10",
X"9d",
X"02",
X"03",
X"a9",
X"04",
X"9d",
X"03",
X"03",
X"a9",
X"00",
X"9d",
X"08",
X"03",
X"8a",
X"18",
X"69",
X"07",
X"8d",
X"00",
X"03",
X"60",
X"ad",
X"33",
X"07",
X"c9",
X"01",
X"d0",
X"05",
X"a9",
X"0b",
X"8d",
X"73",
X"07",
X"4c",
X"45",
X"87",
X"a9",
X"00",
X"20",
X"08",
X"88",
X"4c",
X"45",
X"87",
X"20",
X"30",
X"bc",
X"ae",
X"00",
X"03",
X"a9",
X"20",
X"9d",
X"01",
X"03",
X"a9",
X"73",
X"9d",
X"02",
X"03",
X"a9",
X"03",
X"9d",
X"03",
X"03",
X"ac",
X"5f",
X"07",
X"c8",
X"98",
X"9d",
X"04",
X"03",
X"a9",
X"28",
X"9d",
X"05",
X"03",
X"ac",
X"5c",
X"07",
X"c8",
X"98",
X"9d",
X"06",
X"03",
X"a9",
X"00",
X"9d",
X"07",
X"03",
X"8a",
X"18",
X"69",
X"06",
X"8d",
X"00",
X"03",
X"4c",
X"45",
X"87",
X"ad",
X"59",
X"07",
X"f0",
X"0a",
X"a9",
X"00",
X"8d",
X"59",
X"07",
X"a9",
X"02",
X"4c",
X"c7",
X"86",
X"ee",
X"3c",
X"07",
X"4c",
X"45",
X"87",
X"ad",
X"70",
X"07",
X"f0",
X"33",
X"c9",
X"03",
X"f0",
X"22",
X"ad",
X"52",
X"07",
X"d0",
X"2a",
X"ac",
X"4e",
X"07",
X"c0",
X"03",
X"f0",
X"05",
X"ad",
X"69",
X"07",
X"d0",
X"1e",
X"20",
X"a4",
X"ef",
X"a9",
X"01",
X"20",
X"08",
X"88",
X"20",
X"a5",
X"88",
X"a9",
X"00",
X"8d",
X"74",
X"07",
X"60",
X"a9",
X"12",
X"8d",
X"a0",
X"07",
X"a9",
X"03",
X"20",
X"08",
X"88",
X"4c",
X"4e",
X"87",
X"a9",
X"08",
X"8d",
X"3c",
X"07",
X"60",
X"ee",
X"74",
X"07",
X"20",
X"b0",
X"92",
X"ad",
X"1f",
X"07",
X"d0",
X"f8",
X"ce",
X"1e",
X"07",
X"10",
X"03",
X"ee",
X"3c",
X"07",
X"a9",
X"06",
X"8d",
X"73",
X"07",
X"60",
X"ad",
X"70",
X"07",
X"d0",
X"4a",
X"a9",
X"1e",
X"8d",
X"06",
X"20",
X"a9",
X"c0",
X"8d",
X"06",
X"20",
X"a9",
X"03",
X"85",
X"01",
X"a0",
X"00",
X"84",
X"00",
X"ad",
X"07",
X"20",
X"ad",
X"07",
X"20",
X"91",
X"00",
X"c8",
X"d0",
X"02",
X"e6",
X"01",
X"a5",
X"01",
X"c9",
X"04",
X"d0",
X"f0",
X"c0",
X"3a",
X"90",
X"ec",
X"a9",
X"05",
X"4c",
X"4c",
X"86",
X"ad",
X"70",
X"07",
X"d0",
X"17",
X"a2",
X"00",
X"9d",
X"00",
X"03",
X"9d",
X"00",
X"04",
X"ca",
X"d0",
X"f7",
X"20",
X"25",
X"83",
X"ee",
X"3c",
X"07",
X"60",
X"a9",
X"fa",
X"20",
X"36",
X"bc",
X"ee",
X"72",
X"07",
X"60",
X"20",
X"43",
X"05",
X"16",
X"0a",
X"1b",
X"12",
X"18",
X"20",
X"52",
X"0b",
X"20",
X"18",
X"1b",
X"15",
X"0d",
X"24",
X"24",
X"1d",
X"12",
X"16",
X"0e",
X"20",
X"68",
X"05",
X"00",
X"24",
X"24",
X"2e",
X"29",
X"23",
X"c0",
X"7f",
X"aa",
X"23",
X"c2",
X"01",
X"ea",
X"ff",
X"21",
X"cd",
X"07",
X"24",
X"24",
X"29",
X"24",
X"24",
X"24",
X"24",
X"21",
X"4b",
X"09",
X"20",
X"18",
X"1b",
X"15",
X"0d",
X"24",
X"24",
X"28",
X"24",
X"22",
X"0c",
X"47",
X"24",
X"23",
X"dc",
X"01",
X"ba",
X"ff",
X"21",
X"cd",
X"05",
X"16",
X"0a",
X"1b",
X"12",
X"18",
X"22",
X"0c",
X"07",
X"1d",
X"12",
X"16",
X"0e",
X"24",
X"1e",
X"19",
X"ff",
X"21",
X"cd",
X"05",
X"16",
X"0a",
X"1b",
X"12",
X"18",
X"22",
X"0b",
X"09",
X"10",
X"0a",
X"16",
X"0e",
X"24",
X"18",
X"1f",
X"0e",
X"1b",
X"ff",
X"25",
X"84",
X"15",
X"20",
X"0e",
X"15",
X"0c",
X"18",
X"16",
X"0e",
X"24",
X"1d",
X"18",
X"24",
X"20",
X"0a",
X"1b",
X"19",
X"24",
X"23",
X"18",
X"17",
X"0e",
X"2b",
X"26",
X"25",
X"01",
X"24",
X"26",
X"2d",
X"01",
X"24",
X"26",
X"35",
X"01",
X"24",
X"27",
X"d9",
X"46",
X"aa",
X"27",
X"e1",
X"45",
X"aa",
X"ff",
X"15",
X"1e",
X"12",
X"10",
X"12",
X"04",
X"03",
X"02",
X"00",
X"24",
X"05",
X"24",
X"00",
X"08",
X"07",
X"06",
X"00",
X"00",
X"00",
X"27",
X"27",
X"46",
X"4e",
X"59",
X"61",
X"6e",
X"6e",
X"48",
X"0a",
X"a8",
X"c0",
X"04",
X"90",
X"0c",
X"c0",
X"08",
X"90",
X"02",
X"a0",
X"08",
X"ad",
X"7a",
X"07",
X"d0",
X"01",
X"c8",
X"be",
X"fe",
X"87",
X"a0",
X"00",
X"bd",
X"52",
X"87",
X"c9",
X"ff",
X"f0",
X"07",
X"99",
X"01",
X"03",
X"e8",
X"c8",
X"d0",
X"f2",
X"a9",
X"00",
X"99",
X"01",
X"03",
X"68",
X"aa",
X"c9",
X"04",
X"b0",
X"49",
X"ca",
X"d0",
X"23",
X"ad",
X"5a",
X"07",
X"18",
X"69",
X"01",
X"c9",
X"0a",
X"90",
X"07",
X"e9",
X"0a",
X"a0",
X"9f",
X"8c",
X"08",
X"03",
X"8d",
X"09",
X"03",
X"ac",
X"5f",
X"07",
X"c8",
X"8c",
X"14",
X"03",
X"ac",
X"5c",
X"07",
X"c8",
X"8c",
X"16",
X"03",
X"60",
X"ad",
X"7a",
X"07",
X"f0",
X"1d",
X"ad",
X"53",
X"07",
X"ca",
X"d0",
X"09",
X"ac",
X"70",
X"07",
X"c0",
X"03",
X"f0",
X"02",
X"49",
X"01",
X"4a",
X"90",
X"0b",
X"a0",
X"04",
X"b9",
X"ed",
X"87",
X"99",
X"04",
X"03",
X"88",
X"10",
X"f7",
X"60",
X"e9",
X"04",
X"0a",
X"0a",
X"aa",
X"a0",
X"00",
X"bd",
X"f2",
X"87",
X"99",
X"1c",
X"03",
X"e8",
X"c8",
X"c8",
X"c8",
X"c8",
X"c0",
X"0c",
X"90",
X"f1",
X"a9",
X"2c",
X"4c",
X"3f",
X"86",
X"ad",
X"a0",
X"07",
X"d0",
X"0b",
X"20",
X"20",
X"82",
X"a9",
X"07",
X"8d",
X"a0",
X"07",
X"ee",
X"3c",
X"07",
X"60",
X"ad",
X"26",
X"07",
X"29",
X"01",
X"85",
X"05",
X"ac",
X"40",
X"03",
X"84",
X"00",
X"ad",
X"21",
X"07",
X"99",
X"42",
X"03",
X"ad",
X"20",
X"07",
X"99",
X"41",
X"03",
X"a9",
X"9a",
X"99",
X"43",
X"03",
X"a9",
X"00",
X"85",
X"04",
X"aa",
X"86",
X"01",
X"bd",
X"a1",
X"06",
X"29",
X"c0",
X"85",
X"03",
X"0a",
X"2a",
X"2a",
X"a8",
X"b9",
X"08",
X"8b",
X"85",
X"06",
X"b9",
X"0c",
X"8b",
X"85",
X"07",
X"bd",
X"a1",
X"06",
X"0a",
X"0a",
X"85",
X"02",
X"ad",
X"1f",
X"07",
X"29",
X"01",
X"49",
X"01",
X"0a",
X"65",
X"02",
X"a8",
X"a6",
X"00",
X"b1",
X"06",
X"9d",
X"44",
X"03",
X"c8",
X"b1",
X"06",
X"9d",
X"45",
X"03",
X"a4",
X"04",
X"a5",
X"05",
X"d0",
X"0e",
X"a5",
X"01",
X"4a",
X"b0",
X"19",
X"26",
X"03",
X"26",
X"03",
X"26",
X"03",
X"4c",
X"30",
X"89",
X"a5",
X"01",
X"4a",
X"b0",
X"0f",
X"46",
X"03",
X"46",
X"03",
X"46",
X"03",
X"46",
X"03",
X"4c",
X"30",
X"89",
X"46",
X"03",
X"46",
X"03",
X"e6",
X"04",
X"b9",
X"f9",
X"03",
X"05",
X"03",
X"99",
X"f9",
X"03",
X"e6",
X"00",
X"e6",
X"00",
X"a6",
X"01",
X"e8",
X"e0",
X"0d",
X"90",
X"8d",
X"a4",
X"00",
X"c8",
X"c8",
X"c8",
X"a9",
X"00",
X"99",
X"41",
X"03",
X"8c",
X"40",
X"03",
X"ee",
X"21",
X"07",
X"ad",
X"21",
X"07",
X"29",
X"1f",
X"d0",
X"0d",
X"a9",
X"80",
X"8d",
X"21",
X"07",
X"ad",
X"20",
X"07",
X"49",
X"04",
X"8d",
X"20",
X"07",
X"4c",
X"bd",
X"89",
X"ad",
X"21",
X"07",
X"29",
X"1f",
X"38",
X"e9",
X"04",
X"29",
X"1f",
X"85",
X"01",
X"ad",
X"20",
X"07",
X"b0",
X"02",
X"49",
X"04",
X"29",
X"04",
X"09",
X"23",
X"85",
X"00",
X"a5",
X"01",
X"4a",
X"4a",
X"69",
X"c0",
X"85",
X"01",
X"a2",
X"00",
X"ac",
X"40",
X"03",
X"a5",
X"00",
X"99",
X"41",
X"03",
X"a5",
X"01",
X"18",
X"69",
X"08",
X"99",
X"42",
X"03",
X"85",
X"01",
X"bd",
X"f9",
X"03",
X"99",
X"44",
X"03",
X"a9",
X"01",
X"99",
X"43",
X"03",
X"4a",
X"9d",
X"f9",
X"03",
X"c8",
X"c8",
X"c8",
X"c8",
X"e8",
X"e0",
X"07",
X"90",
X"d9",
X"99",
X"41",
X"03",
X"8c",
X"40",
X"03",
X"a9",
X"06",
X"8d",
X"73",
X"07",
X"60",
X"27",
X"27",
X"27",
X"17",
X"07",
X"17",
X"3f",
X"0c",
X"04",
X"ff",
X"ff",
X"ff",
X"ff",
X"00",
X"0f",
X"07",
X"12",
X"0f",
X"0f",
X"07",
X"17",
X"0f",
X"0f",
X"07",
X"17",
X"1c",
X"0f",
X"07",
X"17",
X"00",
X"a5",
X"09",
X"29",
X"07",
X"d0",
X"51",
X"ae",
X"00",
X"03",
X"e0",
X"31",
X"b0",
X"4a",
X"a8",
X"b9",
X"c9",
X"89",
X"9d",
X"01",
X"03",
X"e8",
X"c8",
X"c0",
X"08",
X"90",
X"f4",
X"ae",
X"00",
X"03",
X"a9",
X"03",
X"85",
X"00",
X"ad",
X"4e",
X"07",
X"0a",
X"0a",
X"a8",
X"b9",
X"d1",
X"89",
X"9d",
X"04",
X"03",
X"c8",
X"e8",
X"c6",
X"00",
X"10",
X"f4",
X"ae",
X"00",
X"03",
X"ac",
X"d4",
X"06",
X"b9",
X"c3",
X"89",
X"9d",
X"05",
X"03",
X"ad",
X"00",
X"03",
X"18",
X"69",
X"07",
X"8d",
X"00",
X"03",
X"ee",
X"d4",
X"06",
X"ad",
X"d4",
X"06",
X"c9",
X"06",
X"90",
X"05",
X"a9",
X"00",
X"8d",
X"d4",
X"06",
X"60",
X"45",
X"45",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"57",
X"58",
X"59",
X"5a",
X"24",
X"24",
X"24",
X"24",
X"26",
X"26",
X"26",
X"26",
X"a0",
X"41",
X"a9",
X"03",
X"ae",
X"4e",
X"07",
X"d0",
X"02",
X"a9",
X"04",
X"20",
X"97",
X"8a",
X"a9",
X"06",
X"8d",
X"73",
X"07",
X"60",
X"20",
X"6d",
X"8a",
X"ee",
X"f0",
X"03",
X"de",
X"ec",
X"03",
X"60",
X"a9",
X"00",
X"a0",
X"03",
X"c9",
X"00",
X"f0",
X"14",
X"a0",
X"00",
X"c9",
X"58",
X"f0",
X"0e",
X"c9",
X"51",
X"f0",
X"0a",
X"c8",
X"c9",
X"5d",
X"f0",
X"05",
X"c9",
X"52",
X"f0",
X"01",
X"c8",
X"98",
X"ac",
X"00",
X"03",
X"c8",
X"20",
X"97",
X"8a",
X"88",
X"98",
X"18",
X"69",
X"0a",
X"4c",
X"3f",
X"86",
X"86",
X"00",
X"84",
X"01",
X"0a",
X"0a",
X"aa",
X"a0",
X"20",
X"a5",
X"06",
X"c9",
X"d0",
X"90",
X"02",
X"a0",
X"24",
X"84",
X"03",
X"29",
X"0f",
X"0a",
X"85",
X"04",
X"a9",
X"00",
X"85",
X"05",
X"a5",
X"02",
X"18",
X"69",
X"20",
X"0a",
X"26",
X"05",
X"0a",
X"26",
X"05",
X"65",
X"04",
X"85",
X"04",
X"a5",
X"05",
X"69",
X"00",
X"18",
X"65",
X"03",
X"85",
X"05",
X"a4",
X"01",
X"bd",
X"39",
X"8a",
X"99",
X"03",
X"03",
X"bd",
X"3a",
X"8a",
X"99",
X"04",
X"03",
X"bd",
X"3b",
X"8a",
X"99",
X"08",
X"03",
X"bd",
X"3c",
X"8a",
X"99",
X"09",
X"03",
X"a5",
X"04",
X"99",
X"01",
X"03",
X"18",
X"69",
X"20",
X"99",
X"06",
X"03",
X"a5",
X"05",
X"99",
X"00",
X"03",
X"99",
X"05",
X"03",
X"a9",
X"02",
X"99",
X"02",
X"03",
X"99",
X"07",
X"03",
X"a9",
X"00",
X"99",
X"0a",
X"03",
X"a6",
X"00",
X"60",
X"10",
X"ac",
X"64",
X"8c",
X"8b",
X"8b",
X"8c",
X"8c",
X"24",
X"24",
X"24",
X"24",
X"27",
X"27",
X"27",
X"27",
X"24",
X"24",
X"24",
X"35",
X"36",
X"25",
X"37",
X"25",
X"24",
X"38",
X"24",
X"24",
X"24",
X"30",
X"30",
X"26",
X"26",
X"26",
X"34",
X"26",
X"24",
X"31",
X"24",
X"32",
X"33",
X"26",
X"24",
X"33",
X"34",
X"26",
X"26",
X"26",
X"26",
X"26",
X"26",
X"26",
X"24",
X"c0",
X"24",
X"c0",
X"24",
X"7f",
X"7f",
X"24",
X"b8",
X"ba",
X"b9",
X"bb",
X"b8",
X"bc",
X"b9",
X"bd",
X"ba",
X"bc",
X"bb",
X"bd",
X"60",
X"64",
X"61",
X"65",
X"62",
X"66",
X"63",
X"67",
X"60",
X"64",
X"61",
X"65",
X"62",
X"66",
X"63",
X"67",
X"68",
X"68",
X"69",
X"69",
X"26",
X"26",
X"6a",
X"6a",
X"4b",
X"4c",
X"4d",
X"4e",
X"4d",
X"4f",
X"4d",
X"4f",
X"4d",
X"4e",
X"50",
X"51",
X"6b",
X"70",
X"2c",
X"2d",
X"6c",
X"71",
X"6d",
X"72",
X"6e",
X"73",
X"6f",
X"74",
X"86",
X"8a",
X"87",
X"8b",
X"88",
X"8c",
X"88",
X"8c",
X"89",
X"8d",
X"69",
X"69",
X"8e",
X"91",
X"8f",
X"92",
X"26",
X"93",
X"26",
X"93",
X"90",
X"94",
X"69",
X"69",
X"a4",
X"e9",
X"ea",
X"eb",
X"24",
X"24",
X"24",
X"24",
X"24",
X"2f",
X"24",
X"3d",
X"a2",
X"a2",
X"a3",
X"a3",
X"24",
X"24",
X"24",
X"24",
X"a2",
X"a2",
X"a3",
X"a3",
X"99",
X"24",
X"99",
X"24",
X"24",
X"a2",
X"3e",
X"3f",
X"5b",
X"5c",
X"24",
X"a3",
X"24",
X"24",
X"24",
X"24",
X"9d",
X"47",
X"9e",
X"47",
X"47",
X"47",
X"27",
X"27",
X"47",
X"47",
X"47",
X"47",
X"27",
X"27",
X"47",
X"47",
X"a9",
X"47",
X"aa",
X"47",
X"9b",
X"27",
X"9c",
X"27",
X"27",
X"27",
X"27",
X"27",
X"52",
X"52",
X"52",
X"52",
X"80",
X"a0",
X"81",
X"a1",
X"be",
X"be",
X"bf",
X"bf",
X"75",
X"ba",
X"76",
X"bb",
X"ba",
X"ba",
X"bb",
X"bb",
X"45",
X"47",
X"45",
X"47",
X"47",
X"47",
X"47",
X"47",
X"45",
X"47",
X"45",
X"47",
X"b4",
X"b6",
X"b5",
X"b7",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"45",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"24",
X"24",
X"24",
X"24",
X"24",
X"24",
X"24",
X"24",
X"ab",
X"ac",
X"ad",
X"ae",
X"5d",
X"5e",
X"5d",
X"5e",
X"c1",
X"24",
X"c1",
X"24",
X"c6",
X"c8",
X"c7",
X"c9",
X"ca",
X"cc",
X"cb",
X"cd",
X"2a",
X"2a",
X"40",
X"40",
X"24",
X"24",
X"24",
X"24",
X"24",
X"47",
X"24",
X"47",
X"82",
X"83",
X"84",
X"85",
X"24",
X"47",
X"24",
X"47",
X"86",
X"8a",
X"87",
X"8b",
X"8e",
X"91",
X"8f",
X"92",
X"24",
X"2f",
X"24",
X"3d",
X"24",
X"24",
X"24",
X"35",
X"36",
X"25",
X"37",
X"25",
X"24",
X"38",
X"24",
X"24",
X"24",
X"24",
X"39",
X"24",
X"3a",
X"24",
X"3b",
X"24",
X"3c",
X"24",
X"24",
X"24",
X"41",
X"26",
X"41",
X"26",
X"26",
X"26",
X"26",
X"26",
X"b0",
X"b1",
X"b2",
X"b3",
X"77",
X"79",
X"77",
X"79",
X"53",
X"55",
X"54",
X"56",
X"53",
X"55",
X"54",
X"56",
X"a5",
X"a7",
X"a6",
X"a8",
X"c2",
X"c4",
X"c3",
X"c5",
X"57",
X"59",
X"58",
X"5a",
X"7b",
X"7d",
X"7c",
X"7e",
X"3f",
X"00",
X"20",
X"0f",
X"15",
X"12",
X"25",
X"0f",
X"3a",
X"1a",
X"0f",
X"0f",
X"30",
X"12",
X"0f",
X"0f",
X"27",
X"12",
X"0f",
X"22",
X"16",
X"27",
X"18",
X"0f",
X"10",
X"30",
X"27",
X"0f",
X"16",
X"30",
X"27",
X"0f",
X"0f",
X"30",
X"10",
X"00",
X"3f",
X"00",
X"20",
X"0f",
X"29",
X"1a",
X"0f",
X"0f",
X"36",
X"17",
X"0f",
X"0f",
X"30",
X"21",
X"0f",
X"0f",
X"27",
X"17",
X"0f",
X"0f",
X"16",
X"27",
X"18",
X"0f",
X"1a",
X"30",
X"27",
X"0f",
X"16",
X"30",
X"27",
X"0f",
X"0f",
X"36",
X"17",
X"00",
X"3f",
X"00",
X"20",
X"0f",
X"29",
X"1a",
X"09",
X"0f",
X"3c",
X"1c",
X"0f",
X"0f",
X"30",
X"21",
X"1c",
X"0f",
X"27",
X"17",
X"1c",
X"0f",
X"16",
X"27",
X"18",
X"0f",
X"1c",
X"36",
X"17",
X"0f",
X"16",
X"30",
X"27",
X"0f",
X"0c",
X"3c",
X"1c",
X"00",
X"3f",
X"00",
X"20",
X"0f",
X"30",
X"10",
X"00",
X"0f",
X"30",
X"10",
X"00",
X"0f",
X"30",
X"16",
X"00",
X"0f",
X"27",
X"17",
X"00",
X"0f",
X"16",
X"27",
X"18",
X"0f",
X"1c",
X"36",
X"17",
X"0f",
X"16",
X"30",
X"27",
X"0f",
X"00",
X"30",
X"10",
X"00",
X"3f",
X"00",
X"04",
X"22",
X"30",
X"00",
X"10",
X"00",
X"3f",
X"00",
X"04",
X"0f",
X"30",
X"00",
X"10",
X"00",
X"3f",
X"00",
X"04",
X"22",
X"27",
X"16",
X"0f",
X"00",
X"3f",
X"14",
X"04",
X"0f",
X"1a",
X"30",
X"27",
X"00",
X"25",
X"48",
X"10",
X"1d",
X"11",
X"0a",
X"17",
X"14",
X"24",
X"22",
X"18",
X"1e",
X"24",
X"16",
X"0a",
X"1b",
X"12",
X"18",
X"2b",
X"00",
X"25",
X"48",
X"10",
X"1d",
X"11",
X"0a",
X"17",
X"14",
X"24",
X"22",
X"18",
X"1e",
X"24",
X"15",
X"1e",
X"12",
X"10",
X"12",
X"2b",
X"00",
X"25",
X"c5",
X"16",
X"0b",
X"1e",
X"1d",
X"24",
X"18",
X"1e",
X"1b",
X"24",
X"19",
X"1b",
X"12",
X"17",
X"0c",
X"0e",
X"1c",
X"1c",
X"24",
X"12",
X"1c",
X"24",
X"12",
X"17",
X"26",
X"05",
X"0f",
X"0a",
X"17",
X"18",
X"1d",
X"11",
X"0e",
X"1b",
X"24",
X"0c",
X"0a",
X"1c",
X"1d",
X"15",
X"0e",
X"2b",
X"00",
X"25",
X"a7",
X"13",
X"22",
X"18",
X"1e",
X"1b",
X"24",
X"1a",
X"1e",
X"0e",
X"1c",
X"1d",
X"24",
X"12",
X"1c",
X"24",
X"18",
X"1f",
X"0e",
X"1b",
X"af",
X"00",
X"25",
X"e3",
X"1b",
X"20",
X"0e",
X"24",
X"19",
X"1b",
X"0e",
X"1c",
X"0e",
X"17",
X"1d",
X"24",
X"22",
X"18",
X"1e",
X"24",
X"0a",
X"24",
X"17",
X"0e",
X"20",
X"24",
X"1a",
X"1e",
X"0e",
X"1c",
X"1d",
X"af",
X"00",
X"26",
X"4a",
X"0d",
X"19",
X"1e",
X"1c",
X"11",
X"24",
X"0b",
X"1e",
X"1d",
X"1d",
X"18",
X"17",
X"24",
X"0b",
X"00",
X"26",
X"88",
X"11",
X"1d",
X"18",
X"24",
X"1c",
X"0e",
X"15",
X"0e",
X"0c",
X"1d",
X"24",
X"0a",
X"24",
X"20",
X"18",
X"1b",
X"15",
X"0d",
X"00",
X"0a",
X"a8",
X"68",
X"85",
X"04",
X"68",
X"85",
X"05",
X"c8",
X"b1",
X"04",
X"85",
X"06",
X"c8",
X"b1",
X"04",
X"85",
X"07",
X"6c",
X"06",
X"00",
X"ad",
X"02",
X"20",
X"ad",
X"78",
X"07",
X"09",
X"10",
X"29",
X"f0",
X"20",
X"ed",
X"8e",
X"a9",
X"24",
X"20",
X"2d",
X"8e",
X"a9",
X"20",
X"8d",
X"06",
X"20",
X"a9",
X"00",
X"8d",
X"06",
X"20",
X"a2",
X"04",
X"a0",
X"c0",
X"a9",
X"24",
X"8d",
X"07",
X"20",
X"88",
X"d0",
X"fa",
X"ca",
X"d0",
X"f7",
X"a0",
X"40",
X"8a",
X"8d",
X"00",
X"03",
X"8d",
X"01",
X"03",
X"8d",
X"07",
X"20",
X"88",
X"d0",
X"fa",
X"8d",
X"3f",
X"07",
X"8d",
X"40",
X"07",
X"4c",
X"e6",
X"8e",
X"a9",
X"01",
X"8d",
X"16",
X"40",
X"4a",
X"aa",
X"8d",
X"16",
X"40",
X"20",
X"6a",
X"8e",
X"e8",
X"a0",
X"08",
X"48",
X"bd",
X"16",
X"40",
X"85",
X"00",
X"4a",
X"05",
X"00",
X"4a",
X"68",
X"2a",
X"88",
X"d0",
X"f1",
X"9d",
X"fc",
X"06",
X"48",
X"29",
X"30",
X"3d",
X"4a",
X"07",
X"f0",
X"07",
X"68",
X"29",
X"cf",
X"9d",
X"fc",
X"06",
X"60",
X"68",
X"9d",
X"4a",
X"07",
X"60",
X"8d",
X"06",
X"20",
X"c8",
X"b1",
X"00",
X"8d",
X"06",
X"20",
X"c8",
X"b1",
X"00",
X"0a",
X"48",
X"ad",
X"78",
X"07",
X"09",
X"04",
X"b0",
X"02",
X"29",
X"fb",
X"20",
X"ed",
X"8e",
X"68",
X"0a",
X"90",
X"03",
X"09",
X"02",
X"c8",
X"4a",
X"4a",
X"aa",
X"b0",
X"01",
X"c8",
X"b1",
X"00",
X"8d",
X"07",
X"20",
X"ca",
X"d0",
X"f5",
X"38",
X"98",
X"65",
X"00",
X"85",
X"00",
X"a9",
X"00",
X"65",
X"01",
X"85",
X"01",
X"a9",
X"3f",
X"8d",
X"06",
X"20",
X"a9",
X"00",
X"8d",
X"06",
X"20",
X"8d",
X"06",
X"20",
X"8d",
X"06",
X"20",
X"ae",
X"02",
X"20",
X"a0",
X"00",
X"b1",
X"00",
X"d0",
X"ac",
X"8d",
X"05",
X"20",
X"8d",
X"05",
X"20",
X"60",
X"8d",
X"00",
X"20",
X"8d",
X"78",
X"07",
X"60",
X"f0",
X"06",
X"62",
X"06",
X"62",
X"06",
X"6d",
X"02",
X"6d",
X"02",
X"7a",
X"03",
X"06",
X"0c",
X"12",
X"18",
X"1e",
X"24",
X"85",
X"00",
X"20",
X"11",
X"8f",
X"a5",
X"00",
X"4a",
X"4a",
X"4a",
X"4a",
X"18",
X"69",
X"01",
X"29",
X"0f",
X"c9",
X"06",
X"b0",
X"44",
X"48",
X"0a",
X"a8",
X"ae",
X"00",
X"03",
X"a9",
X"20",
X"c0",
X"00",
X"d0",
X"02",
X"a9",
X"22",
X"9d",
X"01",
X"03",
X"b9",
X"f4",
X"8e",
X"9d",
X"02",
X"03",
X"b9",
X"f5",
X"8e",
X"9d",
X"03",
X"03",
X"85",
X"03",
X"86",
X"02",
X"68",
X"aa",
X"bd",
X"00",
X"8f",
X"38",
X"f9",
X"f5",
X"8e",
X"a8",
X"a6",
X"02",
X"b9",
X"d7",
X"07",
X"9d",
X"04",
X"03",
X"e8",
X"c8",
X"c6",
X"03",
X"d0",
X"f4",
X"a9",
X"00",
X"9d",
X"04",
X"03",
X"e8",
X"e8",
X"e8",
X"8e",
X"00",
X"03",
X"60",
X"ad",
X"70",
X"07",
X"c9",
X"00",
X"f0",
X"16",
X"a2",
X"05",
X"bd",
X"34",
X"01",
X"18",
X"79",
X"d7",
X"07",
X"30",
X"16",
X"c9",
X"0a",
X"b0",
X"19",
X"99",
X"d7",
X"07",
X"88",
X"ca",
X"10",
X"ec",
X"a9",
X"00",
X"a2",
X"06",
X"9d",
X"33",
X"01",
X"ca",
X"10",
X"fa",
X"60",
X"de",
X"33",
X"01",
X"a9",
X"09",
X"d0",
X"e7",
X"38",
X"e9",
X"0a",
X"fe",
X"33",
X"01",
X"4c",
X"75",
X"8f",
X"a2",
X"05",
X"20",
X"9e",
X"8f",
X"a2",
X"0b",
X"a0",
X"05",
X"38",
X"bd",
X"dd",
X"07",
X"f9",
X"d7",
X"07",
X"ca",
X"88",
X"10",
X"f6",
X"90",
X"0e",
X"e8",
X"c8",
X"bd",
X"dd",
X"07",
X"99",
X"d7",
X"07",
X"e8",
X"c8",
X"c0",
X"06",
X"90",
X"f4",
X"60",
X"04",
X"30",
X"48",
X"60",
X"78",
X"90",
X"a8",
X"c0",
X"d8",
X"e8",
X"24",
X"f8",
X"fc",
X"28",
X"2c",
X"18",
X"ff",
X"23",
X"58",
X"a0",
X"6f",
X"20",
X"cc",
X"90",
X"a0",
X"1f",
X"99",
X"b0",
X"07",
X"88",
X"10",
X"fa",
X"a9",
X"18",
X"8d",
X"a2",
X"07",
X"20",
X"03",
X"9c",
X"a0",
X"4b",
X"20",
X"cc",
X"90",
X"a2",
X"21",
X"a9",
X"00",
X"9d",
X"80",
X"07",
X"ca",
X"10",
X"fa",
X"ad",
X"5b",
X"07",
X"ac",
X"52",
X"07",
X"f0",
X"03",
X"ad",
X"51",
X"07",
X"8d",
X"1a",
X"07",
X"8d",
X"25",
X"07",
X"8d",
X"28",
X"07",
X"20",
X"38",
X"b0",
X"a0",
X"20",
X"29",
X"01",
X"f0",
X"02",
X"a0",
X"24",
X"8c",
X"20",
X"07",
X"a0",
X"80",
X"8c",
X"21",
X"07",
X"0a",
X"0a",
X"0a",
X"0a",
X"8d",
X"a0",
X"06",
X"ce",
X"30",
X"07",
X"ce",
X"31",
X"07",
X"ce",
X"32",
X"07",
X"a9",
X"0b",
X"8d",
X"1e",
X"07",
X"20",
X"22",
X"9c",
X"ad",
X"6a",
X"07",
X"d0",
X"10",
X"ad",
X"5f",
X"07",
X"c9",
X"04",
X"90",
X"0c",
X"d0",
X"07",
X"ad",
X"5c",
X"07",
X"c9",
X"02",
X"90",
X"03",
X"ee",
X"cc",
X"06",
X"ad",
X"5b",
X"07",
X"f0",
X"05",
X"a9",
X"02",
X"8d",
X"10",
X"07",
X"a9",
X"80",
X"85",
X"fb",
X"a9",
X"01",
X"8d",
X"74",
X"07",
X"ee",
X"72",
X"07",
X"60",
X"a9",
X"01",
X"8d",
X"57",
X"07",
X"8d",
X"54",
X"07",
X"a9",
X"02",
X"8d",
X"5a",
X"07",
X"8d",
X"61",
X"07",
X"a9",
X"00",
X"8d",
X"74",
X"07",
X"a8",
X"99",
X"00",
X"03",
X"c8",
X"d0",
X"fa",
X"8d",
X"59",
X"07",
X"8d",
X"69",
X"07",
X"8d",
X"28",
X"07",
X"a9",
X"ff",
X"8d",
X"a0",
X"03",
X"ad",
X"1a",
X"07",
X"4e",
X"78",
X"07",
X"29",
X"01",
X"6a",
X"2e",
X"78",
X"07",
X"20",
X"ed",
X"90",
X"a9",
X"38",
X"8d",
X"e3",
X"06",
X"a9",
X"48",
X"8d",
X"e2",
X"06",
X"a9",
X"58",
X"8d",
X"e1",
X"06",
X"a2",
X"0e",
X"bd",
X"bc",
X"8f",
X"9d",
X"e4",
X"06",
X"ca",
X"10",
X"f7",
X"a0",
X"03",
X"b9",
X"cb",
X"8f",
X"99",
X"00",
X"02",
X"88",
X"10",
X"f7",
X"20",
X"af",
X"92",
X"20",
X"aa",
X"92",
X"ee",
X"22",
X"07",
X"ee",
X"72",
X"07",
X"60",
X"a2",
X"07",
X"a9",
X"00",
X"85",
X"06",
X"86",
X"07",
X"e0",
X"01",
X"d0",
X"04",
X"c0",
X"60",
X"b0",
X"02",
X"91",
X"06",
X"88",
X"c0",
X"ff",
X"d0",
X"f1",
X"ca",
X"10",
X"ec",
X"60",
X"02",
X"01",
X"04",
X"08",
X"10",
X"20",
X"ad",
X"70",
X"07",
X"f0",
X"23",
X"ad",
X"52",
X"07",
X"c9",
X"02",
X"f0",
X"0d",
X"a0",
X"05",
X"ad",
X"10",
X"07",
X"c9",
X"06",
X"f0",
X"0e",
X"c9",
X"07",
X"f0",
X"0a",
X"ac",
X"4e",
X"07",
X"ad",
X"43",
X"07",
X"f0",
X"02",
X"a0",
X"04",
X"b9",
X"e7",
X"90",
X"85",
X"fb",
X"60",
X"28",
X"18",
X"38",
X"28",
X"08",
X"00",
X"00",
X"20",
X"b0",
X"50",
X"00",
X"00",
X"b0",
X"b0",
X"f0",
X"00",
X"20",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"20",
X"04",
X"03",
X"02",
X"ad",
X"1a",
X"07",
X"85",
X"6d",
X"a9",
X"28",
X"8d",
X"0a",
X"07",
X"a9",
X"01",
X"85",
X"33",
X"85",
X"b5",
X"a9",
X"00",
X"85",
X"1d",
X"ce",
X"90",
X"04",
X"a0",
X"00",
X"8c",
X"5b",
X"07",
X"ad",
X"4e",
X"07",
X"d0",
X"01",
X"c8",
X"8c",
X"04",
X"07",
X"ae",
X"10",
X"07",
X"ac",
X"52",
X"07",
X"f0",
X"07",
X"c0",
X"01",
X"f0",
X"03",
X"be",
X"18",
X"91",
X"b9",
X"16",
X"91",
X"85",
X"86",
X"bd",
X"1c",
X"91",
X"85",
X"ce",
X"bd",
X"25",
X"91",
X"8d",
X"c4",
X"03",
X"20",
X"f1",
X"85",
X"ac",
X"15",
X"07",
X"f0",
X"1a",
X"ad",
X"57",
X"07",
X"f0",
X"15",
X"b9",
X"2d",
X"91",
X"8d",
X"f8",
X"07",
X"a9",
X"01",
X"8d",
X"fa",
X"07",
X"4a",
X"8d",
X"f9",
X"07",
X"8d",
X"57",
X"07",
X"8d",
X"9f",
X"07",
X"ac",
X"58",
X"07",
X"f0",
X"14",
X"a9",
X"03",
X"85",
X"1d",
X"a2",
X"00",
X"20",
X"84",
X"bd",
X"a9",
X"f0",
X"85",
X"d7",
X"a2",
X"05",
X"a0",
X"00",
X"20",
X"1e",
X"b9",
X"ac",
X"4e",
X"07",
X"d0",
X"03",
X"20",
X"0b",
X"b7",
X"a9",
X"07",
X"85",
X"0e",
X"60",
X"56",
X"40",
X"65",
X"70",
X"66",
X"40",
X"66",
X"40",
X"66",
X"40",
X"66",
X"60",
X"65",
X"70",
X"00",
X"00",
X"ee",
X"74",
X"07",
X"a9",
X"00",
X"8d",
X"22",
X"07",
X"a9",
X"80",
X"85",
X"fc",
X"ce",
X"5a",
X"07",
X"10",
X"0b",
X"a9",
X"00",
X"8d",
X"72",
X"07",
X"a9",
X"03",
X"8d",
X"70",
X"07",
X"60",
X"ad",
X"5f",
X"07",
X"0a",
X"aa",
X"ad",
X"5c",
X"07",
X"29",
X"02",
X"f0",
X"01",
X"e8",
X"bc",
X"bd",
X"91",
X"ad",
X"5c",
X"07",
X"4a",
X"98",
X"b0",
X"04",
X"4a",
X"4a",
X"4a",
X"4a",
X"29",
X"0f",
X"cd",
X"1a",
X"07",
X"f0",
X"04",
X"90",
X"02",
X"a9",
X"00",
X"8d",
X"5b",
X"07",
X"20",
X"82",
X"92",
X"4c",
X"64",
X"92",
X"ad",
X"72",
X"07",
X"20",
X"04",
X"8e",
X"24",
X"92",
X"67",
X"85",
X"37",
X"92",
X"a9",
X"00",
X"8d",
X"3c",
X"07",
X"8d",
X"22",
X"07",
X"a9",
X"02",
X"85",
X"fc",
X"ee",
X"74",
X"07",
X"ee",
X"72",
X"07",
X"60",
X"a9",
X"00",
X"8d",
X"74",
X"07",
X"ad",
X"fc",
X"06",
X"29",
X"10",
X"d0",
X"05",
X"ad",
X"a0",
X"07",
X"d0",
X"39",
X"a9",
X"80",
X"85",
X"fc",
X"20",
X"82",
X"92",
X"90",
X"13",
X"ad",
X"5f",
X"07",
X"8d",
X"fd",
X"07",
X"a9",
X"00",
X"0a",
X"8d",
X"72",
X"07",
X"8d",
X"a0",
X"07",
X"8d",
X"70",
X"07",
X"60",
X"20",
X"03",
X"9c",
X"a9",
X"01",
X"8d",
X"54",
X"07",
X"ee",
X"57",
X"07",
X"a9",
X"00",
X"8d",
X"47",
X"07",
X"8d",
X"56",
X"07",
X"85",
X"0e",
X"8d",
X"72",
X"07",
X"a9",
X"01",
X"8d",
X"70",
X"07",
X"60",
X"38",
X"ad",
X"7a",
X"07",
X"f0",
X"21",
X"ad",
X"61",
X"07",
X"30",
X"1c",
X"ad",
X"53",
X"07",
X"49",
X"01",
X"8d",
X"53",
X"07",
X"a2",
X"06",
X"bd",
X"5a",
X"07",
X"48",
X"bd",
X"61",
X"07",
X"9d",
X"5a",
X"07",
X"68",
X"9d",
X"61",
X"07",
X"ca",
X"10",
X"ef",
X"18",
X"60",
X"a9",
X"ff",
X"8d",
X"c9",
X"06",
X"60",
X"ac",
X"1f",
X"07",
X"d0",
X"05",
X"a0",
X"08",
X"8c",
X"1f",
X"07",
X"88",
X"98",
X"20",
X"c8",
X"92",
X"ce",
X"1f",
X"07",
X"d0",
X"03",
X"20",
X"6a",
X"89",
X"60",
X"20",
X"04",
X"8e",
X"db",
X"92",
X"ae",
X"88",
X"ae",
X"88",
X"fc",
X"93",
X"db",
X"92",
X"ae",
X"88",
X"ae",
X"88",
X"fc",
X"93",
X"ee",
X"26",
X"07",
X"ad",
X"26",
X"07",
X"29",
X"0f",
X"d0",
X"06",
X"8d",
X"26",
X"07",
X"ee",
X"25",
X"07",
X"ee",
X"a0",
X"06",
X"ad",
X"a0",
X"06",
X"29",
X"1f",
X"8d",
X"a0",
X"06",
X"60",
X"00",
X"30",
X"60",
X"93",
X"00",
X"00",
X"11",
X"12",
X"12",
X"13",
X"00",
X"00",
X"51",
X"52",
X"53",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"91",
X"92",
X"93",
X"00",
X"00",
X"00",
X"00",
X"51",
X"52",
X"53",
X"41",
X"42",
X"43",
X"00",
X"00",
X"00",
X"00",
X"00",
X"91",
X"92",
X"97",
X"87",
X"88",
X"89",
X"99",
X"00",
X"00",
X"00",
X"11",
X"12",
X"13",
X"a4",
X"a5",
X"a5",
X"a5",
X"a6",
X"97",
X"98",
X"99",
X"01",
X"02",
X"03",
X"00",
X"a4",
X"a5",
X"a6",
X"00",
X"11",
X"12",
X"12",
X"12",
X"13",
X"00",
X"00",
X"00",
X"00",
X"01",
X"02",
X"02",
X"03",
X"00",
X"a4",
X"a5",
X"a5",
X"a6",
X"00",
X"00",
X"00",
X"11",
X"12",
X"12",
X"13",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"9c",
X"00",
X"8b",
X"aa",
X"aa",
X"aa",
X"aa",
X"11",
X"12",
X"13",
X"8b",
X"00",
X"9c",
X"9c",
X"00",
X"00",
X"01",
X"02",
X"03",
X"11",
X"12",
X"12",
X"13",
X"00",
X"00",
X"00",
X"00",
X"aa",
X"aa",
X"9c",
X"aa",
X"00",
X"8b",
X"00",
X"01",
X"02",
X"03",
X"80",
X"83",
X"00",
X"81",
X"84",
X"00",
X"82",
X"85",
X"00",
X"02",
X"00",
X"00",
X"03",
X"00",
X"00",
X"04",
X"00",
X"00",
X"00",
X"05",
X"06",
X"07",
X"06",
X"0a",
X"00",
X"08",
X"09",
X"4d",
X"00",
X"00",
X"0d",
X"0f",
X"4e",
X"0e",
X"4e",
X"4e",
X"00",
X"0d",
X"1a",
X"86",
X"87",
X"87",
X"87",
X"87",
X"87",
X"87",
X"87",
X"87",
X"87",
X"87",
X"69",
X"69",
X"00",
X"00",
X"00",
X"00",
X"00",
X"45",
X"47",
X"47",
X"47",
X"47",
X"47",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"86",
X"87",
X"69",
X"54",
X"52",
X"62",
X"00",
X"00",
X"00",
X"18",
X"01",
X"18",
X"07",
X"18",
X"0f",
X"18",
X"ff",
X"18",
X"01",
X"1f",
X"07",
X"1f",
X"0f",
X"1f",
X"81",
X"1f",
X"01",
X"00",
X"8f",
X"1f",
X"f1",
X"1f",
X"f9",
X"18",
X"f1",
X"18",
X"ff",
X"1f",
X"ad",
X"28",
X"07",
X"f0",
X"03",
X"20",
X"08",
X"95",
X"a2",
X"0c",
X"a9",
X"00",
X"9d",
X"a1",
X"06",
X"ca",
X"10",
X"fa",
X"ac",
X"42",
X"07",
X"f0",
X"42",
X"ad",
X"25",
X"07",
X"c9",
X"03",
X"30",
X"05",
X"38",
X"e9",
X"03",
X"10",
X"f7",
X"0a",
X"0a",
X"0a",
X"0a",
X"79",
X"f6",
X"92",
X"6d",
X"26",
X"07",
X"aa",
X"bd",
X"fa",
X"92",
X"f0",
X"26",
X"48",
X"29",
X"0f",
X"38",
X"e9",
X"01",
X"85",
X"00",
X"0a",
X"65",
X"00",
X"aa",
X"68",
X"4a",
X"4a",
X"4a",
X"4a",
X"a8",
X"a9",
X"03",
X"85",
X"00",
X"bd",
X"8a",
X"93",
X"99",
X"a1",
X"06",
X"e8",
X"c8",
X"c0",
X"0b",
X"f0",
X"04",
X"c6",
X"00",
X"d0",
X"f0",
X"ae",
X"41",
X"07",
X"f0",
X"13",
X"bc",
X"ad",
X"93",
X"a2",
X"00",
X"b9",
X"b1",
X"93",
X"f0",
X"03",
X"9d",
X"a1",
X"06",
X"c8",
X"e8",
X"e0",
X"0d",
X"d0",
X"f2",
X"ac",
X"4e",
X"07",
X"d0",
X"0c",
X"ad",
X"5f",
X"07",
X"c9",
X"07",
X"d0",
X"05",
X"a9",
X"62",
X"4c",
X"88",
X"94",
X"b9",
X"d8",
X"93",
X"ac",
X"43",
X"07",
X"f0",
X"02",
X"a9",
X"88",
X"85",
X"07",
X"a2",
X"00",
X"ad",
X"27",
X"07",
X"0a",
X"a8",
X"b9",
X"dc",
X"93",
X"85",
X"00",
X"c8",
X"84",
X"01",
X"ad",
X"43",
X"07",
X"f0",
X"0a",
X"e0",
X"00",
X"f0",
X"06",
X"a5",
X"00",
X"29",
X"08",
X"85",
X"00",
X"a0",
X"00",
X"b9",
X"8a",
X"c6",
X"24",
X"00",
X"f0",
X"05",
X"a5",
X"07",
X"9d",
X"a1",
X"06",
X"e8",
X"e0",
X"0d",
X"f0",
X"18",
X"ad",
X"4e",
X"07",
X"c9",
X"02",
X"d0",
X"08",
X"e0",
X"0b",
X"d0",
X"04",
X"a9",
X"54",
X"85",
X"07",
X"c8",
X"c0",
X"08",
X"d0",
X"db",
X"a4",
X"01",
X"d0",
X"be",
X"20",
X"08",
X"95",
X"ad",
X"a0",
X"06",
X"20",
X"e1",
X"9b",
X"a2",
X"00",
X"a0",
X"00",
X"84",
X"00",
X"bd",
X"a1",
X"06",
X"29",
X"c0",
X"0a",
X"2a",
X"2a",
X"a8",
X"bd",
X"a1",
X"06",
X"d9",
X"04",
X"95",
X"b0",
X"02",
X"a9",
X"00",
X"a4",
X"00",
X"91",
X"06",
X"98",
X"18",
X"69",
X"10",
X"a8",
X"e8",
X"e0",
X"0d",
X"90",
X"dd",
X"60",
X"10",
X"51",
X"88",
X"c0",
X"a2",
X"02",
X"86",
X"08",
X"a9",
X"00",
X"8d",
X"29",
X"07",
X"ac",
X"2c",
X"07",
X"b1",
X"e7",
X"c9",
X"fd",
X"f0",
X"4b",
X"bd",
X"30",
X"07",
X"10",
X"46",
X"c8",
X"b1",
X"e7",
X"0a",
X"90",
X"0b",
X"ad",
X"2b",
X"07",
X"d0",
X"06",
X"ee",
X"2b",
X"07",
X"ee",
X"2a",
X"07",
X"88",
X"b1",
X"e7",
X"29",
X"0f",
X"c9",
X"0d",
X"d0",
X"1b",
X"c8",
X"b1",
X"e7",
X"88",
X"29",
X"40",
X"d0",
X"1c",
X"ad",
X"2b",
X"07",
X"d0",
X"17",
X"c8",
X"b1",
X"e7",
X"29",
X"1f",
X"8d",
X"2a",
X"07",
X"ee",
X"2b",
X"07",
X"4c",
X"6e",
X"95",
X"c9",
X"0e",
X"d0",
X"05",
X"ad",
X"28",
X"07",
X"d0",
X"08",
X"ad",
X"2a",
X"07",
X"cd",
X"25",
X"07",
X"90",
X"06",
X"20",
X"95",
X"95",
X"4c",
X"71",
X"95",
X"ee",
X"29",
X"07",
X"20",
X"89",
X"95",
X"a6",
X"08",
X"bd",
X"30",
X"07",
X"30",
X"03",
X"de",
X"30",
X"07",
X"ca",
X"10",
X"8c",
X"ad",
X"29",
X"07",
X"d0",
X"85",
X"ad",
X"28",
X"07",
X"d0",
X"80",
X"60",
X"ee",
X"2c",
X"07",
X"ee",
X"2c",
X"07",
X"a9",
X"00",
X"8d",
X"2b",
X"07",
X"60",
X"bd",
X"30",
X"07",
X"30",
X"03",
X"bc",
X"2d",
X"07",
X"a2",
X"10",
X"b1",
X"e7",
X"c9",
X"fd",
X"f0",
X"e3",
X"29",
X"0f",
X"c9",
X"0f",
X"f0",
X"08",
X"a2",
X"08",
X"c9",
X"0c",
X"f0",
X"02",
X"a2",
X"00",
X"86",
X"07",
X"a6",
X"08",
X"c9",
X"0e",
X"d0",
X"08",
X"a9",
X"00",
X"85",
X"07",
X"a9",
X"2e",
X"d0",
X"53",
X"c9",
X"0d",
X"d0",
X"1b",
X"a9",
X"22",
X"85",
X"07",
X"c8",
X"b1",
X"e7",
X"29",
X"40",
X"f0",
X"63",
X"b1",
X"e7",
X"29",
X"7f",
X"c9",
X"4b",
X"d0",
X"03",
X"ee",
X"45",
X"07",
X"29",
X"3f",
X"4c",
X"16",
X"96",
X"c9",
X"0c",
X"b0",
X"27",
X"c8",
X"b1",
X"e7",
X"29",
X"70",
X"d0",
X"0b",
X"a9",
X"16",
X"85",
X"07",
X"b1",
X"e7",
X"29",
X"0f",
X"4c",
X"16",
X"96",
X"85",
X"00",
X"c9",
X"70",
X"d0",
X"0a",
X"b1",
X"e7",
X"29",
X"08",
X"f0",
X"04",
X"a9",
X"00",
X"85",
X"00",
X"a5",
X"00",
X"4c",
X"12",
X"96",
X"c8",
X"b1",
X"e7",
X"29",
X"70",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"00",
X"bd",
X"30",
X"07",
X"10",
X"42",
X"ad",
X"2a",
X"07",
X"cd",
X"25",
X"07",
X"f0",
X"11",
X"ac",
X"2c",
X"07",
X"b1",
X"e7",
X"29",
X"0f",
X"c9",
X"0e",
X"d0",
X"05",
X"ad",
X"28",
X"07",
X"d0",
X"21",
X"60",
X"ad",
X"28",
X"07",
X"f0",
X"0b",
X"a9",
X"00",
X"8d",
X"28",
X"07",
X"8d",
X"29",
X"07",
X"85",
X"08",
X"60",
X"ac",
X"2c",
X"07",
X"b1",
X"e7",
X"29",
X"f0",
X"4a",
X"4a",
X"4a",
X"4a",
X"cd",
X"26",
X"07",
X"d0",
X"df",
X"ad",
X"2c",
X"07",
X"9d",
X"2d",
X"07",
X"20",
X"89",
X"95",
X"a5",
X"00",
X"18",
X"65",
X"07",
X"20",
X"04",
X"8e",
X"e5",
X"98",
X"40",
X"97",
X"2e",
X"9a",
X"3e",
X"9a",
X"f2",
X"99",
X"50",
X"9a",
X"59",
X"9a",
X"e5",
X"98",
X"41",
X"9b",
X"ba",
X"97",
X"79",
X"99",
X"7c",
X"99",
X"7f",
X"99",
X"57",
X"99",
X"68",
X"99",
X"6b",
X"99",
X"d0",
X"99",
X"d7",
X"99",
X"06",
X"98",
X"b7",
X"9a",
X"ab",
X"98",
X"94",
X"99",
X"0e",
X"9b",
X"0e",
X"9b",
X"0e",
X"9b",
X"01",
X"9b",
X"19",
X"9b",
X"19",
X"9b",
X"19",
X"9b",
X"14",
X"9b",
X"19",
X"9b",
X"6f",
X"98",
X"19",
X"9a",
X"d3",
X"9a",
X"82",
X"98",
X"9e",
X"99",
X"09",
X"9a",
X"0e",
X"9a",
X"01",
X"9a",
X"f2",
X"96",
X"0d",
X"97",
X"0d",
X"97",
X"2b",
X"97",
X"2b",
X"97",
X"2b",
X"97",
X"45",
X"96",
X"c5",
X"96",
X"bc",
X"2d",
X"07",
X"c8",
X"b1",
X"e7",
X"48",
X"29",
X"40",
X"d0",
X"12",
X"68",
X"48",
X"29",
X"0f",
X"8d",
X"27",
X"07",
X"68",
X"29",
X"30",
X"4a",
X"4a",
X"4a",
X"4a",
X"8d",
X"42",
X"07",
X"60",
X"68",
X"29",
X"07",
X"c9",
X"04",
X"90",
X"05",
X"8d",
X"44",
X"07",
X"a9",
X"00",
X"8d",
X"41",
X"07",
X"60",
X"a2",
X"04",
X"ad",
X"5f",
X"07",
X"f0",
X"08",
X"e8",
X"ac",
X"4e",
X"07",
X"88",
X"d0",
X"01",
X"e8",
X"8a",
X"8d",
X"d6",
X"06",
X"20",
X"08",
X"88",
X"a9",
X"0d",
X"20",
X"16",
X"97",
X"ad",
X"23",
X"07",
X"49",
X"01",
X"8d",
X"23",
X"07",
X"60",
X"85",
X"00",
X"a9",
X"00",
X"a2",
X"04",
X"b4",
X"16",
X"c4",
X"00",
X"d0",
X"02",
X"95",
X"0f",
X"ca",
X"10",
X"f5",
X"60",
X"14",
X"17",
X"18",
X"a6",
X"00",
X"bd",
X"20",
X"97",
X"a0",
X"05",
X"88",
X"30",
X"07",
X"d9",
X"16",
X"00",
X"d0",
X"f8",
X"a9",
X"00",
X"8d",
X"cd",
X"06",
X"60",
X"ad",
X"33",
X"07",
X"20",
X"04",
X"8e",
X"4c",
X"97",
X"78",
X"97",
X"69",
X"9a",
X"20",
X"bb",
X"9b",
X"bd",
X"30",
X"07",
X"f0",
X"1f",
X"10",
X"11",
X"98",
X"9d",
X"30",
X"07",
X"ad",
X"25",
X"07",
X"0d",
X"26",
X"07",
X"f0",
X"05",
X"a9",
X"16",
X"4c",
X"b0",
X"97",
X"a6",
X"07",
X"a9",
X"17",
X"9d",
X"a1",
X"06",
X"a9",
X"4c",
X"4c",
X"aa",
X"97",
X"a9",
X"18",
X"4c",
X"b0",
X"97",
X"20",
X"ac",
X"9b",
X"84",
X"06",
X"90",
X"0c",
X"bd",
X"30",
X"07",
X"4a",
X"9d",
X"36",
X"07",
X"a9",
X"19",
X"4c",
X"b0",
X"97",
X"a9",
X"1b",
X"bc",
X"30",
X"07",
X"f0",
X"1e",
X"bd",
X"36",
X"07",
X"85",
X"06",
X"a6",
X"07",
X"a9",
X"1a",
X"9d",
X"a1",
X"06",
X"c4",
X"06",
X"d0",
X"2c",
X"e8",
X"a9",
X"4f",
X"9d",
X"a1",
X"06",
X"a9",
X"50",
X"e8",
X"a0",
X"0f",
X"4c",
X"7d",
X"9b",
X"a6",
X"07",
X"a0",
X"00",
X"4c",
X"7d",
X"9b",
X"42",
X"41",
X"43",
X"20",
X"ac",
X"9b",
X"a0",
X"00",
X"b0",
X"07",
X"c8",
X"bd",
X"30",
X"07",
X"d0",
X"01",
X"c8",
X"b9",
X"b7",
X"97",
X"8d",
X"a1",
X"06",
X"60",
X"00",
X"45",
X"45",
X"45",
X"00",
X"00",
X"48",
X"47",
X"46",
X"00",
X"45",
X"49",
X"49",
X"49",
X"45",
X"47",
X"47",
X"4a",
X"47",
X"47",
X"47",
X"47",
X"4b",
X"47",
X"47",
X"49",
X"49",
X"49",
X"49",
X"49",
X"47",
X"4a",
X"47",
X"4a",
X"47",
X"47",
X"4b",
X"47",
X"4b",
X"47",
X"47",
X"47",
X"47",
X"47",
X"47",
X"4a",
X"47",
X"4a",
X"47",
X"4a",
X"4b",
X"47",
X"4b",
X"47",
X"4b",
X"20",
X"bb",
X"9b",
X"84",
X"07",
X"a0",
X"04",
X"20",
X"af",
X"9b",
X"8a",
X"48",
X"bc",
X"30",
X"07",
X"a6",
X"07",
X"a9",
X"0b",
X"85",
X"06",
X"b9",
X"cf",
X"97",
X"9d",
X"a1",
X"06",
X"e8",
X"a5",
X"06",
X"f0",
X"07",
X"c8",
X"c8",
X"c8",
X"c8",
X"c8",
X"c6",
X"06",
X"e0",
X"0b",
X"d0",
X"ea",
X"68",
X"aa",
X"ad",
X"25",
X"07",
X"f0",
X"36",
X"bd",
X"30",
X"07",
X"c9",
X"01",
X"f0",
X"2a",
X"a4",
X"07",
X"d0",
X"04",
X"c9",
X"03",
X"f0",
X"22",
X"c9",
X"02",
X"d0",
X"23",
X"20",
X"cb",
X"9b",
X"48",
X"20",
X"4a",
X"99",
X"68",
X"95",
X"87",
X"ad",
X"25",
X"07",
X"95",
X"6e",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"a9",
X"90",
X"95",
X"cf",
X"a9",
X"31",
X"95",
X"16",
X"60",
X"a0",
X"52",
X"8c",
X"ab",
X"06",
X"60",
X"20",
X"bb",
X"9b",
X"bc",
X"30",
X"07",
X"a6",
X"07",
X"a9",
X"6b",
X"9d",
X"a1",
X"06",
X"a9",
X"6c",
X"9d",
X"a2",
X"06",
X"60",
X"a0",
X"03",
X"20",
X"af",
X"9b",
X"a0",
X"0a",
X"20",
X"b3",
X"98",
X"b0",
X"10",
X"a2",
X"06",
X"a9",
X"00",
X"9d",
X"a1",
X"06",
X"ca",
X"10",
X"f8",
X"b9",
X"dd",
X"98",
X"8d",
X"a8",
X"06",
X"60",
X"15",
X"14",
X"00",
X"00",
X"15",
X"1e",
X"1d",
X"1c",
X"15",
X"21",
X"20",
X"1f",
X"a0",
X"03",
X"20",
X"af",
X"9b",
X"20",
X"bb",
X"9b",
X"88",
X"88",
X"84",
X"05",
X"bc",
X"30",
X"07",
X"84",
X"06",
X"a6",
X"05",
X"e8",
X"b9",
X"9f",
X"98",
X"c9",
X"00",
X"f0",
X"08",
X"a2",
X"00",
X"a4",
X"05",
X"20",
X"7d",
X"9b",
X"18",
X"a4",
X"06",
X"b9",
X"a3",
X"98",
X"9d",
X"a1",
X"06",
X"b9",
X"a7",
X"98",
X"9d",
X"a2",
X"06",
X"60",
X"11",
X"10",
X"15",
X"14",
X"13",
X"12",
X"15",
X"14",
X"20",
X"39",
X"99",
X"a5",
X"00",
X"f0",
X"04",
X"c8",
X"c8",
X"c8",
X"c8",
X"98",
X"48",
X"ad",
X"60",
X"07",
X"0d",
X"5f",
X"07",
X"f0",
X"2b",
X"bc",
X"30",
X"07",
X"f0",
X"26",
X"20",
X"4a",
X"99",
X"b0",
X"21",
X"20",
X"cb",
X"9b",
X"18",
X"69",
X"08",
X"95",
X"87",
X"ad",
X"25",
X"07",
X"69",
X"00",
X"95",
X"6e",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"20",
X"d3",
X"9b",
X"95",
X"cf",
X"a9",
X"0d",
X"95",
X"16",
X"20",
X"87",
X"c7",
X"68",
X"a8",
X"a6",
X"07",
X"b9",
X"dd",
X"98",
X"9d",
X"a1",
X"06",
X"e8",
X"b9",
X"df",
X"98",
X"a4",
X"06",
X"88",
X"4c",
X"7d",
X"9b",
X"a0",
X"01",
X"20",
X"af",
X"9b",
X"20",
X"bb",
X"9b",
X"98",
X"29",
X"07",
X"85",
X"06",
X"bc",
X"30",
X"07",
X"60",
X"a2",
X"00",
X"18",
X"b5",
X"0f",
X"f0",
X"05",
X"e8",
X"e0",
X"05",
X"d0",
X"f6",
X"60",
X"20",
X"ac",
X"9b",
X"a9",
X"86",
X"8d",
X"ab",
X"06",
X"a2",
X"0b",
X"a0",
X"01",
X"a9",
X"87",
X"4c",
X"7d",
X"9b",
X"a9",
X"03",
X"2c",
X"a9",
X"07",
X"48",
X"20",
X"ac",
X"9b",
X"68",
X"aa",
X"a9",
X"c0",
X"9d",
X"a1",
X"06",
X"60",
X"a9",
X"06",
X"2c",
X"a9",
X"07",
X"2c",
X"a9",
X"09",
X"48",
X"20",
X"ac",
X"9b",
X"68",
X"aa",
X"a9",
X"0b",
X"9d",
X"a1",
X"06",
X"e8",
X"a0",
X"00",
X"a9",
X"63",
X"4c",
X"7d",
X"9b",
X"20",
X"bb",
X"9b",
X"a2",
X"02",
X"a9",
X"6d",
X"4c",
X"7d",
X"9b",
X"a9",
X"24",
X"8d",
X"a1",
X"06",
X"a2",
X"01",
X"a0",
X"08",
X"a9",
X"25",
X"20",
X"7d",
X"9b",
X"a9",
X"61",
X"8d",
X"ab",
X"06",
X"20",
X"cb",
X"9b",
X"38",
X"e9",
X"08",
X"85",
X"8c",
X"ad",
X"25",
X"07",
X"e9",
X"00",
X"85",
X"73",
X"a9",
X"30",
X"85",
X"d4",
X"a9",
X"b0",
X"8d",
X"0d",
X"01",
X"a9",
X"30",
X"85",
X"1b",
X"e6",
X"14",
X"60",
X"a2",
X"00",
X"a0",
X"0f",
X"4c",
X"e9",
X"99",
X"8a",
X"48",
X"a2",
X"01",
X"a0",
X"0f",
X"a9",
X"44",
X"20",
X"7d",
X"9b",
X"68",
X"aa",
X"20",
X"bb",
X"9b",
X"a2",
X"01",
X"a9",
X"40",
X"4c",
X"7d",
X"9b",
X"c3",
X"c2",
X"c2",
X"c2",
X"ac",
X"4e",
X"07",
X"b9",
X"ee",
X"99",
X"4c",
X"44",
X"9a",
X"06",
X"07",
X"08",
X"c5",
X"0c",
X"89",
X"a0",
X"0c",
X"20",
X"af",
X"9b",
X"4c",
X"0e",
X"9a",
X"a9",
X"08",
X"8d",
X"73",
X"07",
X"a4",
X"00",
X"be",
X"f9",
X"99",
X"b9",
X"fc",
X"99",
X"4c",
X"20",
X"9a",
X"20",
X"bb",
X"9b",
X"a6",
X"07",
X"a9",
X"c4",
X"a0",
X"00",
X"4c",
X"7d",
X"9b",
X"69",
X"61",
X"61",
X"62",
X"22",
X"51",
X"52",
X"52",
X"88",
X"ac",
X"4e",
X"07",
X"ad",
X"43",
X"07",
X"f0",
X"02",
X"a0",
X"04",
X"b9",
X"29",
X"9a",
X"4c",
X"44",
X"9a",
X"ac",
X"4e",
X"07",
X"b9",
X"25",
X"9a",
X"48",
X"20",
X"ac",
X"9b",
X"a6",
X"07",
X"a0",
X"00",
X"68",
X"4c",
X"7d",
X"9b",
X"ac",
X"4e",
X"07",
X"b9",
X"29",
X"9a",
X"4c",
X"5f",
X"9a",
X"ac",
X"4e",
X"07",
X"b9",
X"25",
X"9a",
X"48",
X"20",
X"bb",
X"9b",
X"68",
X"a6",
X"07",
X"4c",
X"7d",
X"9b",
X"20",
X"bb",
X"9b",
X"a6",
X"07",
X"a9",
X"64",
X"9d",
X"a1",
X"06",
X"e8",
X"88",
X"30",
X"0e",
X"a9",
X"65",
X"9d",
X"a1",
X"06",
X"e8",
X"88",
X"30",
X"05",
X"a9",
X"66",
X"20",
X"7d",
X"9b",
X"ae",
X"6a",
X"04",
X"20",
X"d3",
X"9b",
X"9d",
X"77",
X"04",
X"ad",
X"25",
X"07",
X"9d",
X"6b",
X"04",
X"20",
X"cb",
X"9b",
X"9d",
X"71",
X"04",
X"e8",
X"e0",
X"06",
X"90",
X"02",
X"a2",
X"00",
X"8e",
X"6a",
X"04",
X"60",
X"07",
X"07",
X"06",
X"05",
X"04",
X"03",
X"02",
X"01",
X"00",
X"03",
X"03",
X"04",
X"05",
X"06",
X"07",
X"08",
X"09",
X"0a",
X"20",
X"ac",
X"9b",
X"90",
X"05",
X"a9",
X"09",
X"8d",
X"34",
X"07",
X"ce",
X"34",
X"07",
X"ac",
X"34",
X"07",
X"be",
X"ae",
X"9a",
X"b9",
X"a5",
X"9a",
X"a8",
X"a9",
X"61",
X"4c",
X"7d",
X"9b",
X"20",
X"bb",
X"9b",
X"20",
X"4a",
X"99",
X"20",
X"cb",
X"9b",
X"95",
X"87",
X"ad",
X"25",
X"07",
X"95",
X"6e",
X"20",
X"d3",
X"9b",
X"95",
X"cf",
X"95",
X"58",
X"a9",
X"32",
X"95",
X"16",
X"a0",
X"01",
X"94",
X"b6",
X"f6",
X"0f",
X"a6",
X"07",
X"a9",
X"67",
X"9d",
X"a1",
X"06",
X"a9",
X"68",
X"9d",
X"a2",
X"06",
X"60",
X"ad",
X"5d",
X"07",
X"f0",
X"36",
X"a9",
X"00",
X"8d",
X"5d",
X"07",
X"4c",
X"19",
X"9b",
X"20",
X"36",
X"9b",
X"4c",
X"2c",
X"9b",
X"a9",
X"00",
X"8d",
X"bc",
X"06",
X"20",
X"36",
X"9b",
X"84",
X"07",
X"a9",
X"00",
X"ac",
X"4e",
X"07",
X"88",
X"f0",
X"02",
X"a9",
X"05",
X"18",
X"65",
X"07",
X"a8",
X"b9",
X"e8",
X"bd",
X"48",
X"20",
X"bb",
X"9b",
X"4c",
X"48",
X"9a",
X"a5",
X"00",
X"38",
X"e9",
X"00",
X"a8",
X"60",
X"87",
X"00",
X"00",
X"00",
X"20",
X"ac",
X"9b",
X"90",
X"2d",
X"ad",
X"4e",
X"07",
X"d0",
X"28",
X"ae",
X"6a",
X"04",
X"20",
X"cb",
X"9b",
X"38",
X"e9",
X"10",
X"9d",
X"71",
X"04",
X"ad",
X"25",
X"07",
X"e9",
X"00",
X"9d",
X"6b",
X"04",
X"c8",
X"c8",
X"98",
X"0a",
X"0a",
X"0a",
X"0a",
X"9d",
X"77",
X"04",
X"e8",
X"e0",
X"05",
X"90",
X"02",
X"a2",
X"00",
X"8e",
X"6a",
X"04",
X"ae",
X"4e",
X"07",
X"bd",
X"3d",
X"9b",
X"a2",
X"08",
X"a0",
X"0f",
X"8c",
X"35",
X"07",
X"bc",
X"a1",
X"06",
X"f0",
X"18",
X"c0",
X"17",
X"f0",
X"17",
X"c0",
X"1a",
X"f0",
X"13",
X"c0",
X"c0",
X"f0",
X"0c",
X"c0",
X"c0",
X"b0",
X"0b",
X"c0",
X"54",
X"d0",
X"04",
X"c9",
X"50",
X"f0",
X"03",
X"9d",
X"a1",
X"06",
X"e8",
X"e0",
X"0d",
X"b0",
X"06",
X"ac",
X"35",
X"07",
X"88",
X"10",
X"d2",
X"60",
X"20",
X"bb",
X"9b",
X"bd",
X"30",
X"07",
X"18",
X"10",
X"05",
X"98",
X"9d",
X"30",
X"07",
X"38",
X"60",
X"bc",
X"2d",
X"07",
X"b1",
X"e7",
X"29",
X"0f",
X"85",
X"07",
X"c8",
X"b1",
X"e7",
X"29",
X"0f",
X"a8",
X"60",
X"ad",
X"26",
X"07",
X"0a",
X"0a",
X"0a",
X"0a",
X"60",
X"a5",
X"07",
X"0a",
X"0a",
X"0a",
X"0a",
X"18",
X"69",
X"20",
X"60",
X"00",
X"d0",
X"05",
X"05",
X"48",
X"4a",
X"4a",
X"4a",
X"4a",
X"a8",
X"b9",
X"df",
X"9b",
X"85",
X"07",
X"68",
X"29",
X"0f",
X"18",
X"79",
X"dd",
X"9b",
X"85",
X"06",
X"60",
X"ff",
X"ff",
X"12",
X"36",
X"0e",
X"0e",
X"0e",
X"32",
X"32",
X"32",
X"0a",
X"26",
X"40",
X"20",
X"13",
X"9c",
X"8d",
X"50",
X"07",
X"29",
X"60",
X"0a",
X"2a",
X"2a",
X"2a",
X"8d",
X"4e",
X"07",
X"60",
X"ac",
X"5f",
X"07",
X"b9",
X"b4",
X"9c",
X"18",
X"6d",
X"60",
X"07",
X"a8",
X"b9",
X"bc",
X"9c",
X"60",
X"ad",
X"50",
X"07",
X"20",
X"09",
X"9c",
X"a8",
X"ad",
X"50",
X"07",
X"29",
X"1f",
X"8d",
X"4f",
X"07",
X"b9",
X"e0",
X"9c",
X"18",
X"6d",
X"4f",
X"07",
X"a8",
X"b9",
X"e4",
X"9c",
X"85",
X"e9",
X"b9",
X"06",
X"9d",
X"85",
X"ea",
X"ac",
X"4e",
X"07",
X"b9",
X"28",
X"9d",
X"18",
X"6d",
X"4f",
X"07",
X"a8",
X"b9",
X"2c",
X"9d",
X"85",
X"e7",
X"b9",
X"4e",
X"9d",
X"85",
X"e8",
X"a0",
X"00",
X"b1",
X"e7",
X"48",
X"29",
X"07",
X"c9",
X"04",
X"90",
X"05",
X"8d",
X"44",
X"07",
X"a9",
X"00",
X"8d",
X"41",
X"07",
X"68",
X"48",
X"29",
X"38",
X"4a",
X"4a",
X"4a",
X"8d",
X"10",
X"07",
X"68",
X"29",
X"c0",
X"18",
X"2a",
X"2a",
X"2a",
X"8d",
X"15",
X"07",
X"c8",
X"b1",
X"e7",
X"48",
X"29",
X"0f",
X"8d",
X"27",
X"07",
X"68",
X"48",
X"29",
X"30",
X"4a",
X"4a",
X"4a",
X"4a",
X"8d",
X"42",
X"07",
X"68",
X"29",
X"c0",
X"18",
X"2a",
X"2a",
X"2a",
X"c9",
X"03",
X"d0",
X"05",
X"8d",
X"43",
X"07",
X"a9",
X"00",
X"8d",
X"33",
X"07",
X"a5",
X"e7",
X"18",
X"69",
X"02",
X"85",
X"e7",
X"a5",
X"e8",
X"69",
X"00",
X"85",
X"e8",
X"60",
X"00",
X"05",
X"0a",
X"0e",
X"13",
X"17",
X"1b",
X"20",
X"25",
X"29",
X"c0",
X"26",
X"60",
X"28",
X"29",
X"01",
X"27",
X"62",
X"24",
X"35",
X"20",
X"63",
X"22",
X"29",
X"41",
X"2c",
X"61",
X"2a",
X"31",
X"26",
X"62",
X"2e",
X"23",
X"2d",
X"60",
X"33",
X"29",
X"01",
X"27",
X"64",
X"30",
X"32",
X"21",
X"65",
X"1f",
X"06",
X"1c",
X"00",
X"70",
X"97",
X"b0",
X"df",
X"0a",
X"1f",
X"59",
X"7e",
X"9b",
X"a9",
X"d0",
X"01",
X"1f",
X"3c",
X"51",
X"7b",
X"7c",
X"a0",
X"a9",
X"ce",
X"f1",
X"fa",
X"fb",
X"35",
X"60",
X"8e",
X"aa",
X"b3",
X"d8",
X"05",
X"33",
X"60",
X"71",
X"9b",
X"9d",
X"9d",
X"9d",
X"9d",
X"9e",
X"9e",
X"9e",
X"9e",
X"9e",
X"9e",
X"9e",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"9f",
X"a0",
X"a0",
X"a0",
X"a0",
X"a0",
X"a0",
X"a1",
X"a1",
X"a1",
X"a1",
X"a1",
X"00",
X"03",
X"19",
X"1c",
X"06",
X"45",
X"c0",
X"6b",
X"ce",
X"37",
X"8a",
X"19",
X"8e",
X"f3",
X"48",
X"cd",
X"32",
X"3b",
X"7a",
X"8f",
X"f6",
X"5b",
X"ce",
X"ff",
X"92",
X"05",
X"7e",
X"d7",
X"02",
X"35",
X"d8",
X"79",
X"af",
X"10",
X"8f",
X"02",
X"6f",
X"fa",
X"ae",
X"ae",
X"ae",
X"a4",
X"a4",
X"a5",
X"a5",
X"a6",
X"a6",
X"a6",
X"a7",
X"a7",
X"a8",
X"a8",
X"a8",
X"a8",
X"a8",
X"a9",
X"a9",
X"a9",
X"aa",
X"ab",
X"ab",
X"ab",
X"ac",
X"ac",
X"ac",
X"ad",
X"a1",
X"a2",
X"a2",
X"a3",
X"a3",
X"a3",
X"76",
X"dd",
X"bb",
X"4c",
X"ea",
X"1d",
X"1b",
X"cc",
X"56",
X"5d",
X"16",
X"9d",
X"c6",
X"1d",
X"36",
X"9d",
X"c9",
X"1d",
X"04",
X"db",
X"49",
X"1d",
X"84",
X"1b",
X"c9",
X"5d",
X"88",
X"95",
X"0f",
X"08",
X"30",
X"4c",
X"78",
X"2d",
X"a6",
X"28",
X"90",
X"b5",
X"ff",
X"0f",
X"03",
X"56",
X"1b",
X"c9",
X"1b",
X"0f",
X"07",
X"36",
X"1b",
X"aa",
X"1b",
X"48",
X"95",
X"0f",
X"0a",
X"2a",
X"1b",
X"5b",
X"0c",
X"78",
X"2d",
X"90",
X"b5",
X"ff",
X"0b",
X"8c",
X"4b",
X"4c",
X"77",
X"5f",
X"eb",
X"0c",
X"bd",
X"db",
X"19",
X"9d",
X"75",
X"1d",
X"7d",
X"5b",
X"d9",
X"1d",
X"3d",
X"dd",
X"99",
X"1d",
X"26",
X"9d",
X"5a",
X"2b",
X"8a",
X"2c",
X"ca",
X"1b",
X"20",
X"95",
X"7b",
X"5c",
X"db",
X"4c",
X"1b",
X"cc",
X"3b",
X"cc",
X"78",
X"2d",
X"a6",
X"28",
X"90",
X"b5",
X"ff",
X"0b",
X"8c",
X"3b",
X"1d",
X"8b",
X"1d",
X"ab",
X"0c",
X"db",
X"1d",
X"0f",
X"03",
X"65",
X"1d",
X"6b",
X"1b",
X"05",
X"9d",
X"0b",
X"1b",
X"05",
X"9b",
X"0b",
X"1d",
X"8b",
X"0c",
X"1b",
X"8c",
X"70",
X"15",
X"7b",
X"0c",
X"db",
X"0c",
X"0f",
X"08",
X"78",
X"2d",
X"a6",
X"28",
X"90",
X"b5",
X"ff",
X"27",
X"a9",
X"4b",
X"0c",
X"68",
X"29",
X"0f",
X"06",
X"77",
X"1b",
X"0f",
X"0b",
X"60",
X"15",
X"4b",
X"8c",
X"78",
X"2d",
X"90",
X"b5",
X"ff",
X"0f",
X"03",
X"8e",
X"65",
X"e1",
X"bb",
X"38",
X"6d",
X"a8",
X"3e",
X"e5",
X"e7",
X"0f",
X"08",
X"0b",
X"02",
X"2b",
X"02",
X"5e",
X"65",
X"e1",
X"bb",
X"0e",
X"db",
X"0e",
X"bb",
X"8e",
X"db",
X"0e",
X"fe",
X"65",
X"ec",
X"0f",
X"0d",
X"4e",
X"65",
X"e1",
X"0f",
X"0e",
X"4e",
X"02",
X"e0",
X"0f",
X"10",
X"fe",
X"e5",
X"e1",
X"1b",
X"85",
X"7b",
X"0c",
X"5b",
X"95",
X"78",
X"2d",
X"90",
X"b5",
X"ff",
X"a5",
X"86",
X"e4",
X"28",
X"18",
X"a8",
X"45",
X"83",
X"69",
X"03",
X"c6",
X"29",
X"9b",
X"83",
X"16",
X"a4",
X"88",
X"24",
X"e9",
X"28",
X"05",
X"a8",
X"7b",
X"28",
X"24",
X"8f",
X"c8",
X"03",
X"e8",
X"03",
X"46",
X"a8",
X"85",
X"24",
X"c8",
X"24",
X"ff",
X"eb",
X"8e",
X"0f",
X"03",
X"fb",
X"05",
X"17",
X"85",
X"db",
X"8e",
X"0f",
X"07",
X"57",
X"05",
X"7b",
X"05",
X"9b",
X"80",
X"2b",
X"85",
X"fb",
X"05",
X"0f",
X"0b",
X"1b",
X"05",
X"9b",
X"05",
X"ff",
X"2e",
X"c2",
X"66",
X"e2",
X"11",
X"0f",
X"07",
X"02",
X"11",
X"0f",
X"0c",
X"12",
X"11",
X"ff",
X"0e",
X"c2",
X"a8",
X"ab",
X"00",
X"bb",
X"8e",
X"6b",
X"82",
X"de",
X"00",
X"a0",
X"33",
X"86",
X"43",
X"06",
X"3e",
X"b4",
X"a0",
X"cb",
X"02",
X"0f",
X"07",
X"7e",
X"42",
X"a6",
X"83",
X"02",
X"0f",
X"0a",
X"3b",
X"02",
X"cb",
X"37",
X"0f",
X"0c",
X"e3",
X"0e",
X"ff",
X"9b",
X"8e",
X"ca",
X"0e",
X"ee",
X"42",
X"44",
X"5b",
X"86",
X"80",
X"b8",
X"1b",
X"80",
X"50",
X"ba",
X"10",
X"b7",
X"5b",
X"00",
X"17",
X"85",
X"4b",
X"05",
X"fe",
X"34",
X"40",
X"b7",
X"86",
X"c6",
X"06",
X"5b",
X"80",
X"83",
X"00",
X"d0",
X"38",
X"5b",
X"8e",
X"8a",
X"0e",
X"a6",
X"00",
X"bb",
X"0e",
X"c5",
X"80",
X"f3",
X"00",
X"ff",
X"1e",
X"c2",
X"00",
X"6b",
X"06",
X"8b",
X"86",
X"63",
X"b7",
X"0f",
X"05",
X"03",
X"06",
X"23",
X"06",
X"4b",
X"b7",
X"bb",
X"00",
X"5b",
X"b7",
X"fb",
X"37",
X"3b",
X"b7",
X"0f",
X"0b",
X"1b",
X"37",
X"ff",
X"2b",
X"d7",
X"e3",
X"03",
X"c2",
X"86",
X"e2",
X"06",
X"76",
X"a5",
X"a3",
X"8f",
X"03",
X"86",
X"2b",
X"57",
X"68",
X"28",
X"e9",
X"28",
X"e5",
X"83",
X"24",
X"8f",
X"36",
X"a8",
X"5b",
X"03",
X"ff",
X"0f",
X"02",
X"78",
X"40",
X"48",
X"ce",
X"f8",
X"c3",
X"f8",
X"c3",
X"0f",
X"07",
X"7b",
X"43",
X"c6",
X"d0",
X"0f",
X"8a",
X"c8",
X"50",
X"ff",
X"85",
X"86",
X"0b",
X"80",
X"1b",
X"00",
X"db",
X"37",
X"77",
X"80",
X"eb",
X"37",
X"fe",
X"2b",
X"20",
X"2b",
X"80",
X"7b",
X"38",
X"ab",
X"b8",
X"77",
X"86",
X"fe",
X"42",
X"20",
X"49",
X"86",
X"8b",
X"06",
X"9b",
X"80",
X"7b",
X"8e",
X"5b",
X"b7",
X"9b",
X"0e",
X"bb",
X"0e",
X"9b",
X"80",
X"ff",
X"0b",
X"80",
X"60",
X"38",
X"10",
X"b8",
X"c0",
X"3b",
X"db",
X"8e",
X"40",
X"b8",
X"f0",
X"38",
X"7b",
X"8e",
X"a0",
X"b8",
X"c0",
X"b8",
X"fb",
X"00",
X"a0",
X"b8",
X"30",
X"bb",
X"ee",
X"42",
X"88",
X"0f",
X"0b",
X"2b",
X"0e",
X"67",
X"0e",
X"ff",
X"0a",
X"aa",
X"0e",
X"28",
X"2a",
X"0e",
X"31",
X"88",
X"ff",
X"c7",
X"83",
X"d7",
X"03",
X"42",
X"8f",
X"7a",
X"03",
X"05",
X"a4",
X"78",
X"24",
X"a6",
X"25",
X"e4",
X"25",
X"4b",
X"83",
X"e3",
X"03",
X"05",
X"a4",
X"89",
X"24",
X"b5",
X"24",
X"09",
X"a4",
X"65",
X"24",
X"c9",
X"24",
X"0f",
X"08",
X"85",
X"25",
X"ff",
X"cd",
X"a5",
X"b5",
X"a8",
X"07",
X"a8",
X"76",
X"28",
X"cc",
X"25",
X"65",
X"a4",
X"a9",
X"24",
X"e5",
X"24",
X"19",
X"a4",
X"0f",
X"07",
X"95",
X"28",
X"e6",
X"24",
X"19",
X"a4",
X"d7",
X"29",
X"16",
X"a9",
X"58",
X"29",
X"97",
X"29",
X"ff",
X"0f",
X"02",
X"02",
X"11",
X"0f",
X"07",
X"02",
X"11",
X"ff",
X"ff",
X"2b",
X"82",
X"ab",
X"38",
X"de",
X"42",
X"e2",
X"1b",
X"b8",
X"eb",
X"3b",
X"db",
X"80",
X"8b",
X"b8",
X"1b",
X"82",
X"fb",
X"b8",
X"7b",
X"80",
X"fb",
X"3c",
X"5b",
X"bc",
X"7b",
X"b8",
X"1b",
X"8e",
X"cb",
X"0e",
X"1b",
X"8e",
X"0f",
X"0d",
X"2b",
X"3b",
X"bb",
X"b8",
X"eb",
X"82",
X"4b",
X"b8",
X"bb",
X"38",
X"3b",
X"b7",
X"bb",
X"02",
X"0f",
X"13",
X"1b",
X"00",
X"cb",
X"80",
X"6b",
X"bc",
X"ff",
X"7b",
X"80",
X"ae",
X"00",
X"80",
X"8b",
X"8e",
X"e8",
X"05",
X"f9",
X"86",
X"17",
X"86",
X"16",
X"85",
X"4e",
X"2b",
X"80",
X"ab",
X"8e",
X"87",
X"85",
X"c3",
X"05",
X"8b",
X"82",
X"9b",
X"02",
X"ab",
X"02",
X"bb",
X"86",
X"cb",
X"06",
X"d3",
X"03",
X"3b",
X"8e",
X"6b",
X"0e",
X"a7",
X"8e",
X"ff",
X"29",
X"8e",
X"52",
X"11",
X"83",
X"0e",
X"0f",
X"03",
X"9b",
X"0e",
X"2b",
X"8e",
X"5b",
X"0e",
X"cb",
X"8e",
X"fb",
X"0e",
X"fb",
X"82",
X"9b",
X"82",
X"bb",
X"02",
X"fe",
X"42",
X"e8",
X"bb",
X"8e",
X"0f",
X"0a",
X"ab",
X"0e",
X"cb",
X"0e",
X"f9",
X"0e",
X"88",
X"86",
X"a6",
X"06",
X"db",
X"02",
X"b6",
X"8e",
X"ff",
X"ab",
X"ce",
X"de",
X"42",
X"c0",
X"cb",
X"ce",
X"5b",
X"8e",
X"1b",
X"ce",
X"4b",
X"85",
X"67",
X"45",
X"0f",
X"07",
X"2b",
X"00",
X"7b",
X"85",
X"97",
X"05",
X"0f",
X"0a",
X"92",
X"02",
X"ff",
X"0a",
X"aa",
X"0e",
X"24",
X"4a",
X"1e",
X"23",
X"aa",
X"ff",
X"1b",
X"80",
X"bb",
X"38",
X"4b",
X"bc",
X"eb",
X"3b",
X"0f",
X"04",
X"2b",
X"00",
X"ab",
X"38",
X"eb",
X"00",
X"cb",
X"8e",
X"fb",
X"80",
X"ab",
X"b8",
X"6b",
X"80",
X"fb",
X"3c",
X"9b",
X"bb",
X"5b",
X"bc",
X"fb",
X"00",
X"6b",
X"b8",
X"fb",
X"38",
X"ff",
X"0b",
X"86",
X"1a",
X"06",
X"db",
X"06",
X"de",
X"c2",
X"02",
X"f0",
X"3b",
X"bb",
X"80",
X"eb",
X"06",
X"0b",
X"86",
X"93",
X"06",
X"f0",
X"39",
X"0f",
X"06",
X"60",
X"b8",
X"1b",
X"86",
X"a0",
X"b9",
X"b7",
X"27",
X"bd",
X"27",
X"2b",
X"83",
X"a1",
X"26",
X"a9",
X"26",
X"ee",
X"25",
X"0b",
X"27",
X"b4",
X"ff",
X"0f",
X"02",
X"1e",
X"2f",
X"60",
X"e0",
X"3a",
X"a5",
X"a7",
X"db",
X"80",
X"3b",
X"82",
X"8b",
X"02",
X"fe",
X"42",
X"68",
X"70",
X"bb",
X"25",
X"a7",
X"2c",
X"27",
X"b2",
X"26",
X"b9",
X"26",
X"9b",
X"80",
X"a8",
X"82",
X"b5",
X"27",
X"bc",
X"27",
X"b0",
X"bb",
X"3b",
X"82",
X"87",
X"34",
X"ee",
X"25",
X"6b",
X"ff",
X"1e",
X"a5",
X"0a",
X"2e",
X"28",
X"27",
X"2e",
X"33",
X"c7",
X"0f",
X"03",
X"1e",
X"40",
X"07",
X"2e",
X"30",
X"e7",
X"0f",
X"05",
X"1e",
X"24",
X"44",
X"0f",
X"07",
X"1e",
X"22",
X"6a",
X"2e",
X"23",
X"ab",
X"0f",
X"09",
X"1e",
X"41",
X"68",
X"1e",
X"2a",
X"8a",
X"2e",
X"23",
X"a2",
X"2e",
X"32",
X"ea",
X"ff",
X"3b",
X"87",
X"66",
X"27",
X"cc",
X"27",
X"ee",
X"31",
X"87",
X"ee",
X"23",
X"a7",
X"3b",
X"87",
X"db",
X"07",
X"ff",
X"0f",
X"01",
X"2e",
X"25",
X"2b",
X"2e",
X"25",
X"4b",
X"4e",
X"25",
X"cb",
X"6b",
X"07",
X"97",
X"47",
X"e9",
X"87",
X"47",
X"c7",
X"7a",
X"07",
X"d6",
X"c7",
X"78",
X"07",
X"38",
X"87",
X"ab",
X"47",
X"e3",
X"07",
X"9b",
X"87",
X"0f",
X"09",
X"68",
X"47",
X"db",
X"c7",
X"3b",
X"c7",
X"ff",
X"47",
X"9b",
X"cb",
X"07",
X"fa",
X"1d",
X"86",
X"9b",
X"3a",
X"87",
X"56",
X"07",
X"88",
X"1b",
X"07",
X"9d",
X"2e",
X"65",
X"f0",
X"ff",
X"9b",
X"07",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"ce",
X"03",
X"dc",
X"51",
X"ee",
X"07",
X"73",
X"e0",
X"74",
X"0a",
X"7e",
X"06",
X"9e",
X"0a",
X"ce",
X"06",
X"e4",
X"00",
X"e8",
X"0a",
X"fe",
X"0a",
X"2e",
X"89",
X"4e",
X"0b",
X"54",
X"0a",
X"14",
X"8a",
X"c4",
X"0a",
X"34",
X"8a",
X"7e",
X"06",
X"c7",
X"0a",
X"01",
X"e0",
X"02",
X"0a",
X"47",
X"0a",
X"81",
X"60",
X"82",
X"0a",
X"c7",
X"0a",
X"0e",
X"87",
X"7e",
X"02",
X"a7",
X"02",
X"b3",
X"02",
X"d7",
X"02",
X"e3",
X"02",
X"07",
X"82",
X"13",
X"02",
X"3e",
X"06",
X"7e",
X"02",
X"ae",
X"07",
X"fe",
X"0a",
X"0d",
X"c4",
X"cd",
X"43",
X"ce",
X"09",
X"de",
X"0b",
X"dd",
X"42",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"5b",
X"07",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"5e",
X"0a",
X"68",
X"64",
X"98",
X"64",
X"a8",
X"64",
X"ce",
X"06",
X"fe",
X"02",
X"0d",
X"01",
X"1e",
X"0e",
X"7e",
X"02",
X"94",
X"63",
X"b4",
X"63",
X"d4",
X"63",
X"f4",
X"63",
X"14",
X"e3",
X"2e",
X"0e",
X"5e",
X"02",
X"64",
X"35",
X"88",
X"72",
X"be",
X"0e",
X"0d",
X"04",
X"ae",
X"02",
X"ce",
X"08",
X"cd",
X"4b",
X"fe",
X"02",
X"0d",
X"05",
X"68",
X"31",
X"7e",
X"0a",
X"96",
X"31",
X"a9",
X"63",
X"a8",
X"33",
X"d5",
X"30",
X"ee",
X"02",
X"e6",
X"62",
X"f4",
X"61",
X"04",
X"b1",
X"08",
X"3f",
X"44",
X"33",
X"94",
X"63",
X"a4",
X"31",
X"e4",
X"31",
X"04",
X"bf",
X"08",
X"3f",
X"04",
X"bf",
X"08",
X"3f",
X"cd",
X"4b",
X"03",
X"e4",
X"0e",
X"03",
X"2e",
X"01",
X"7e",
X"06",
X"be",
X"02",
X"de",
X"06",
X"fe",
X"0a",
X"0d",
X"c4",
X"cd",
X"43",
X"ce",
X"09",
X"de",
X"0b",
X"dd",
X"42",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"9b",
X"07",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"fe",
X"00",
X"27",
X"b1",
X"65",
X"32",
X"75",
X"0a",
X"71",
X"00",
X"b7",
X"31",
X"08",
X"e4",
X"18",
X"64",
X"1e",
X"04",
X"57",
X"3b",
X"bb",
X"0a",
X"17",
X"8a",
X"27",
X"3a",
X"73",
X"0a",
X"7b",
X"0a",
X"d7",
X"0a",
X"e7",
X"3a",
X"3b",
X"8a",
X"97",
X"0a",
X"fe",
X"08",
X"24",
X"8a",
X"2e",
X"00",
X"3e",
X"40",
X"38",
X"64",
X"6f",
X"00",
X"9f",
X"00",
X"be",
X"43",
X"c8",
X"0a",
X"c9",
X"63",
X"ce",
X"07",
X"fe",
X"07",
X"2e",
X"81",
X"66",
X"42",
X"6a",
X"42",
X"79",
X"0a",
X"be",
X"00",
X"c8",
X"64",
X"f8",
X"64",
X"08",
X"e4",
X"2e",
X"07",
X"7e",
X"03",
X"9e",
X"07",
X"be",
X"03",
X"de",
X"07",
X"fe",
X"0a",
X"03",
X"a5",
X"0d",
X"44",
X"cd",
X"43",
X"ce",
X"09",
X"dd",
X"42",
X"de",
X"0b",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"9b",
X"07",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"fe",
X"06",
X"0c",
X"81",
X"39",
X"0a",
X"5c",
X"01",
X"89",
X"0a",
X"ac",
X"01",
X"d9",
X"0a",
X"fc",
X"01",
X"2e",
X"83",
X"a7",
X"01",
X"b7",
X"00",
X"c7",
X"01",
X"de",
X"0a",
X"fe",
X"02",
X"4e",
X"83",
X"5a",
X"32",
X"63",
X"0a",
X"69",
X"0a",
X"7e",
X"02",
X"ee",
X"03",
X"fa",
X"32",
X"03",
X"8a",
X"09",
X"0a",
X"1e",
X"02",
X"ee",
X"03",
X"fa",
X"32",
X"03",
X"8a",
X"09",
X"0a",
X"14",
X"42",
X"1e",
X"02",
X"7e",
X"0a",
X"9e",
X"07",
X"fe",
X"0a",
X"2e",
X"86",
X"5e",
X"0a",
X"8e",
X"06",
X"be",
X"0a",
X"ee",
X"07",
X"3e",
X"83",
X"5e",
X"07",
X"fe",
X"0a",
X"0d",
X"c4",
X"41",
X"52",
X"51",
X"52",
X"cd",
X"43",
X"ce",
X"09",
X"de",
X"0b",
X"dd",
X"42",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"5b",
X"07",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"fe",
X"0a",
X"ae",
X"86",
X"be",
X"07",
X"fe",
X"02",
X"0d",
X"02",
X"27",
X"32",
X"46",
X"61",
X"55",
X"62",
X"5e",
X"0e",
X"1e",
X"82",
X"68",
X"3c",
X"74",
X"3a",
X"7d",
X"4b",
X"5e",
X"8e",
X"7d",
X"4b",
X"7e",
X"82",
X"84",
X"62",
X"94",
X"61",
X"a4",
X"31",
X"bd",
X"4b",
X"ce",
X"06",
X"fe",
X"02",
X"0d",
X"06",
X"34",
X"31",
X"3e",
X"0a",
X"64",
X"32",
X"75",
X"0a",
X"7b",
X"61",
X"a4",
X"33",
X"ae",
X"02",
X"de",
X"0e",
X"3e",
X"82",
X"64",
X"32",
X"78",
X"32",
X"b4",
X"36",
X"c8",
X"36",
X"dd",
X"4b",
X"44",
X"b2",
X"58",
X"32",
X"94",
X"63",
X"a4",
X"3e",
X"ba",
X"30",
X"c9",
X"61",
X"ce",
X"06",
X"dd",
X"4b",
X"ce",
X"86",
X"dd",
X"4b",
X"fe",
X"02",
X"2e",
X"86",
X"5e",
X"02",
X"7e",
X"06",
X"fe",
X"02",
X"1e",
X"86",
X"3e",
X"02",
X"5e",
X"06",
X"7e",
X"02",
X"9e",
X"06",
X"fe",
X"0a",
X"0d",
X"c4",
X"cd",
X"43",
X"ce",
X"09",
X"de",
X"0b",
X"dd",
X"42",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"5b",
X"06",
X"05",
X"32",
X"06",
X"33",
X"07",
X"34",
X"5e",
X"0a",
X"ae",
X"02",
X"0d",
X"01",
X"39",
X"73",
X"0d",
X"03",
X"39",
X"7b",
X"4d",
X"4b",
X"de",
X"06",
X"1e",
X"8a",
X"ae",
X"06",
X"c4",
X"33",
X"16",
X"fe",
X"a5",
X"77",
X"fe",
X"02",
X"fe",
X"82",
X"0d",
X"07",
X"39",
X"73",
X"a8",
X"74",
X"ed",
X"4b",
X"49",
X"fb",
X"e8",
X"74",
X"fe",
X"0a",
X"2e",
X"82",
X"67",
X"02",
X"84",
X"7a",
X"87",
X"31",
X"0d",
X"0b",
X"fe",
X"02",
X"0d",
X"0c",
X"39",
X"73",
X"5e",
X"06",
X"c6",
X"76",
X"45",
X"ff",
X"be",
X"0a",
X"dd",
X"48",
X"fe",
X"06",
X"3d",
X"cb",
X"46",
X"7e",
X"ad",
X"4a",
X"fe",
X"82",
X"39",
X"f3",
X"a9",
X"7b",
X"4e",
X"8a",
X"9e",
X"07",
X"fe",
X"0a",
X"0d",
X"c4",
X"cd",
X"43",
X"ce",
X"09",
X"de",
X"0b",
X"dd",
X"42",
X"fe",
X"02",
X"5d",
X"c7",
X"fd",
X"94",
X"11",
X"0f",
X"26",
X"fe",
X"10",
X"28",
X"94",
X"65",
X"15",
X"eb",
X"12",
X"fa",
X"41",
X"4a",
X"96",
X"54",
X"40",
X"a4",
X"42",
X"b7",
X"13",
X"e9",
X"19",
X"f5",
X"15",
X"11",
X"80",
X"47",
X"42",
X"71",
X"13",
X"80",
X"41",
X"15",
X"92",
X"1b",
X"1f",
X"24",
X"40",
X"55",
X"12",
X"64",
X"40",
X"95",
X"12",
X"a4",
X"40",
X"d2",
X"12",
X"e1",
X"40",
X"13",
X"c0",
X"2c",
X"17",
X"2f",
X"12",
X"49",
X"13",
X"83",
X"40",
X"9f",
X"14",
X"a3",
X"40",
X"17",
X"92",
X"83",
X"13",
X"92",
X"41",
X"b9",
X"14",
X"c5",
X"12",
X"c8",
X"40",
X"d4",
X"40",
X"4b",
X"92",
X"78",
X"1b",
X"9c",
X"94",
X"9f",
X"11",
X"df",
X"14",
X"fe",
X"11",
X"7d",
X"c1",
X"9e",
X"42",
X"cf",
X"20",
X"fd",
X"90",
X"b1",
X"0f",
X"26",
X"29",
X"91",
X"7e",
X"42",
X"fe",
X"40",
X"28",
X"92",
X"4e",
X"42",
X"2e",
X"c0",
X"57",
X"73",
X"c3",
X"25",
X"c7",
X"27",
X"23",
X"84",
X"33",
X"20",
X"5c",
X"01",
X"77",
X"63",
X"88",
X"62",
X"99",
X"61",
X"aa",
X"60",
X"bc",
X"01",
X"ee",
X"42",
X"4e",
X"c0",
X"69",
X"11",
X"7e",
X"42",
X"de",
X"40",
X"f8",
X"62",
X"0e",
X"c2",
X"ae",
X"40",
X"d7",
X"63",
X"e7",
X"63",
X"33",
X"a7",
X"37",
X"27",
X"43",
X"04",
X"cc",
X"01",
X"e7",
X"73",
X"0c",
X"81",
X"3e",
X"42",
X"0d",
X"0a",
X"5e",
X"40",
X"88",
X"72",
X"be",
X"42",
X"e7",
X"87",
X"fe",
X"40",
X"39",
X"e1",
X"4e",
X"00",
X"69",
X"60",
X"87",
X"60",
X"a5",
X"60",
X"c3",
X"31",
X"fe",
X"31",
X"6d",
X"c1",
X"be",
X"42",
X"ef",
X"20",
X"fd",
X"52",
X"21",
X"0f",
X"20",
X"6e",
X"40",
X"58",
X"f2",
X"93",
X"01",
X"97",
X"00",
X"0c",
X"81",
X"97",
X"40",
X"a6",
X"41",
X"c7",
X"40",
X"0d",
X"04",
X"03",
X"01",
X"07",
X"01",
X"23",
X"01",
X"27",
X"01",
X"ec",
X"03",
X"ac",
X"f3",
X"c3",
X"03",
X"78",
X"e2",
X"94",
X"43",
X"47",
X"f3",
X"74",
X"43",
X"47",
X"fb",
X"74",
X"43",
X"2c",
X"f1",
X"4c",
X"63",
X"47",
X"00",
X"57",
X"21",
X"5c",
X"01",
X"7c",
X"72",
X"39",
X"f1",
X"ec",
X"02",
X"4c",
X"81",
X"d8",
X"62",
X"ec",
X"01",
X"0d",
X"0d",
X"0f",
X"38",
X"c7",
X"07",
X"ed",
X"4a",
X"1d",
X"c1",
X"5f",
X"26",
X"fd",
X"54",
X"21",
X"0f",
X"26",
X"a7",
X"22",
X"37",
X"fb",
X"73",
X"20",
X"83",
X"07",
X"87",
X"02",
X"93",
X"20",
X"c7",
X"73",
X"04",
X"f1",
X"06",
X"31",
X"39",
X"71",
X"59",
X"71",
X"e7",
X"73",
X"37",
X"a0",
X"47",
X"04",
X"86",
X"7c",
X"e5",
X"71",
X"e7",
X"31",
X"33",
X"a4",
X"39",
X"71",
X"a9",
X"71",
X"d3",
X"23",
X"08",
X"f2",
X"13",
X"05",
X"27",
X"02",
X"49",
X"71",
X"75",
X"75",
X"e8",
X"72",
X"67",
X"f3",
X"99",
X"71",
X"e7",
X"20",
X"f4",
X"72",
X"f7",
X"31",
X"17",
X"a0",
X"33",
X"20",
X"39",
X"71",
X"73",
X"28",
X"bc",
X"05",
X"39",
X"f1",
X"79",
X"71",
X"a6",
X"21",
X"c3",
X"06",
X"d3",
X"20",
X"dc",
X"00",
X"fc",
X"00",
X"07",
X"a2",
X"13",
X"21",
X"5f",
X"32",
X"8c",
X"00",
X"98",
X"7a",
X"c7",
X"63",
X"d9",
X"61",
X"03",
X"a2",
X"07",
X"22",
X"74",
X"72",
X"77",
X"31",
X"e7",
X"73",
X"39",
X"f1",
X"58",
X"72",
X"77",
X"73",
X"d8",
X"72",
X"7f",
X"b1",
X"97",
X"73",
X"b6",
X"64",
X"c5",
X"65",
X"d4",
X"66",
X"e3",
X"67",
X"f3",
X"67",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"52",
X"31",
X"0f",
X"20",
X"6e",
X"66",
X"07",
X"81",
X"36",
X"01",
X"66",
X"00",
X"a7",
X"22",
X"08",
X"f2",
X"67",
X"7b",
X"dc",
X"02",
X"98",
X"f2",
X"d7",
X"20",
X"39",
X"f1",
X"9f",
X"33",
X"dc",
X"27",
X"dc",
X"57",
X"23",
X"83",
X"57",
X"63",
X"6c",
X"51",
X"87",
X"63",
X"99",
X"61",
X"a3",
X"06",
X"b3",
X"21",
X"77",
X"f3",
X"f3",
X"21",
X"f7",
X"2a",
X"13",
X"81",
X"23",
X"22",
X"53",
X"00",
X"63",
X"22",
X"e9",
X"0b",
X"0c",
X"83",
X"13",
X"21",
X"16",
X"22",
X"33",
X"05",
X"8f",
X"35",
X"ec",
X"01",
X"63",
X"a0",
X"67",
X"20",
X"73",
X"01",
X"77",
X"01",
X"83",
X"20",
X"87",
X"20",
X"b3",
X"20",
X"b7",
X"20",
X"c3",
X"01",
X"c7",
X"00",
X"d3",
X"20",
X"d7",
X"20",
X"67",
X"a0",
X"77",
X"07",
X"87",
X"22",
X"e8",
X"62",
X"f5",
X"65",
X"1c",
X"82",
X"7f",
X"38",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"50",
X"21",
X"07",
X"81",
X"47",
X"24",
X"57",
X"00",
X"63",
X"01",
X"77",
X"01",
X"c9",
X"71",
X"68",
X"f2",
X"e7",
X"73",
X"97",
X"fb",
X"06",
X"83",
X"5c",
X"01",
X"d7",
X"22",
X"e7",
X"00",
X"03",
X"a7",
X"6c",
X"02",
X"b3",
X"22",
X"e3",
X"01",
X"e7",
X"07",
X"47",
X"a0",
X"57",
X"06",
X"a7",
X"01",
X"d3",
X"00",
X"d7",
X"01",
X"07",
X"81",
X"67",
X"20",
X"93",
X"22",
X"03",
X"a3",
X"1c",
X"61",
X"17",
X"21",
X"6f",
X"33",
X"c7",
X"63",
X"d8",
X"62",
X"e9",
X"61",
X"fa",
X"60",
X"4f",
X"b3",
X"87",
X"63",
X"9c",
X"01",
X"b7",
X"63",
X"c8",
X"62",
X"d9",
X"61",
X"ea",
X"60",
X"39",
X"f1",
X"87",
X"21",
X"a7",
X"01",
X"b7",
X"20",
X"39",
X"f1",
X"5f",
X"38",
X"6d",
X"c1",
X"af",
X"26",
X"fd",
X"90",
X"11",
X"0f",
X"26",
X"fe",
X"10",
X"2a",
X"93",
X"87",
X"17",
X"a3",
X"14",
X"b2",
X"42",
X"0a",
X"92",
X"19",
X"40",
X"36",
X"14",
X"50",
X"41",
X"82",
X"16",
X"2b",
X"93",
X"24",
X"41",
X"bb",
X"14",
X"b8",
X"00",
X"c2",
X"43",
X"c3",
X"13",
X"1b",
X"94",
X"67",
X"12",
X"c4",
X"15",
X"53",
X"c1",
X"d2",
X"41",
X"12",
X"c1",
X"29",
X"13",
X"85",
X"17",
X"1b",
X"92",
X"1a",
X"42",
X"47",
X"13",
X"83",
X"41",
X"a7",
X"13",
X"0e",
X"91",
X"a7",
X"63",
X"b7",
X"63",
X"c5",
X"65",
X"d5",
X"65",
X"dd",
X"4a",
X"e3",
X"67",
X"f3",
X"67",
X"8d",
X"c1",
X"ae",
X"42",
X"df",
X"20",
X"fd",
X"90",
X"11",
X"0f",
X"26",
X"6e",
X"10",
X"8b",
X"17",
X"af",
X"32",
X"d8",
X"62",
X"e8",
X"62",
X"fc",
X"3f",
X"ad",
X"c8",
X"f8",
X"64",
X"0c",
X"be",
X"43",
X"43",
X"f8",
X"64",
X"0c",
X"bf",
X"73",
X"40",
X"84",
X"40",
X"93",
X"40",
X"a4",
X"40",
X"b3",
X"40",
X"f8",
X"64",
X"48",
X"e4",
X"5c",
X"39",
X"83",
X"40",
X"92",
X"41",
X"b3",
X"40",
X"f8",
X"64",
X"48",
X"e4",
X"5c",
X"39",
X"f8",
X"64",
X"13",
X"c2",
X"37",
X"65",
X"4c",
X"24",
X"63",
X"00",
X"97",
X"65",
X"c3",
X"42",
X"0b",
X"97",
X"ac",
X"32",
X"f8",
X"64",
X"0c",
X"be",
X"53",
X"45",
X"9d",
X"48",
X"f8",
X"64",
X"2a",
X"e2",
X"3c",
X"47",
X"56",
X"43",
X"ba",
X"62",
X"f8",
X"64",
X"0c",
X"b7",
X"88",
X"64",
X"bc",
X"31",
X"d4",
X"45",
X"fc",
X"31",
X"3c",
X"b1",
X"78",
X"64",
X"8c",
X"38",
X"0b",
X"9c",
X"1a",
X"33",
X"18",
X"61",
X"28",
X"61",
X"39",
X"60",
X"5d",
X"4a",
X"ee",
X"11",
X"0f",
X"b8",
X"1d",
X"c1",
X"3e",
X"42",
X"6f",
X"20",
X"fd",
X"52",
X"31",
X"0f",
X"20",
X"6e",
X"40",
X"f7",
X"20",
X"07",
X"84",
X"17",
X"20",
X"4f",
X"34",
X"c3",
X"03",
X"c7",
X"02",
X"d3",
X"22",
X"27",
X"e3",
X"39",
X"61",
X"e7",
X"73",
X"5c",
X"e4",
X"57",
X"00",
X"6c",
X"73",
X"47",
X"a0",
X"53",
X"06",
X"63",
X"22",
X"a7",
X"73",
X"fc",
X"73",
X"13",
X"a1",
X"33",
X"05",
X"43",
X"21",
X"5c",
X"72",
X"c3",
X"23",
X"cc",
X"03",
X"77",
X"fb",
X"ac",
X"02",
X"39",
X"f1",
X"a7",
X"73",
X"d3",
X"04",
X"e8",
X"72",
X"e3",
X"22",
X"26",
X"f4",
X"bc",
X"02",
X"8c",
X"81",
X"a8",
X"62",
X"17",
X"87",
X"43",
X"24",
X"a7",
X"01",
X"c3",
X"04",
X"08",
X"f2",
X"97",
X"21",
X"a3",
X"02",
X"c9",
X"0b",
X"e1",
X"69",
X"f1",
X"69",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"38",
X"11",
X"0f",
X"26",
X"ad",
X"40",
X"3d",
X"c7",
X"fd",
X"95",
X"b1",
X"0f",
X"26",
X"0d",
X"02",
X"c8",
X"72",
X"1c",
X"81",
X"38",
X"72",
X"0d",
X"05",
X"97",
X"34",
X"98",
X"62",
X"a3",
X"20",
X"b3",
X"06",
X"c3",
X"20",
X"cc",
X"03",
X"f9",
X"91",
X"2c",
X"81",
X"48",
X"62",
X"0d",
X"09",
X"37",
X"63",
X"47",
X"03",
X"57",
X"21",
X"8c",
X"02",
X"c5",
X"79",
X"c7",
X"31",
X"f9",
X"11",
X"39",
X"f1",
X"a9",
X"11",
X"6f",
X"b4",
X"d3",
X"65",
X"e3",
X"65",
X"7d",
X"c1",
X"bf",
X"26",
X"fd",
X"00",
X"c1",
X"4c",
X"00",
X"f4",
X"4f",
X"0d",
X"02",
X"02",
X"42",
X"43",
X"4f",
X"52",
X"c2",
X"de",
X"00",
X"5a",
X"c2",
X"4d",
X"c7",
X"fd",
X"90",
X"51",
X"0f",
X"26",
X"ee",
X"10",
X"0b",
X"94",
X"33",
X"14",
X"42",
X"42",
X"77",
X"16",
X"86",
X"44",
X"02",
X"92",
X"4a",
X"16",
X"69",
X"42",
X"73",
X"14",
X"b0",
X"00",
X"c7",
X"12",
X"05",
X"c0",
X"1c",
X"17",
X"1f",
X"11",
X"36",
X"12",
X"8f",
X"14",
X"91",
X"40",
X"1b",
X"94",
X"35",
X"12",
X"34",
X"42",
X"60",
X"42",
X"61",
X"12",
X"87",
X"12",
X"96",
X"40",
X"a3",
X"14",
X"1c",
X"98",
X"1f",
X"11",
X"47",
X"12",
X"9f",
X"15",
X"cc",
X"15",
X"cf",
X"11",
X"05",
X"c0",
X"1f",
X"15",
X"39",
X"12",
X"7c",
X"16",
X"7f",
X"11",
X"82",
X"40",
X"98",
X"12",
X"df",
X"15",
X"16",
X"c4",
X"17",
X"14",
X"54",
X"12",
X"9b",
X"16",
X"28",
X"94",
X"ce",
X"01",
X"3d",
X"c1",
X"5e",
X"42",
X"8f",
X"20",
X"fd",
X"97",
X"11",
X"0f",
X"26",
X"fe",
X"10",
X"2b",
X"92",
X"57",
X"12",
X"8b",
X"12",
X"c0",
X"41",
X"f7",
X"13",
X"5b",
X"92",
X"69",
X"0b",
X"bb",
X"12",
X"b2",
X"46",
X"19",
X"93",
X"71",
X"00",
X"17",
X"94",
X"7c",
X"14",
X"7f",
X"11",
X"93",
X"41",
X"bf",
X"15",
X"fc",
X"13",
X"ff",
X"11",
X"2f",
X"95",
X"50",
X"42",
X"51",
X"12",
X"58",
X"14",
X"a6",
X"12",
X"db",
X"12",
X"1b",
X"93",
X"46",
X"43",
X"7b",
X"12",
X"8d",
X"49",
X"b7",
X"14",
X"1b",
X"94",
X"49",
X"0b",
X"bb",
X"12",
X"fc",
X"13",
X"ff",
X"12",
X"03",
X"c1",
X"2f",
X"15",
X"43",
X"12",
X"4b",
X"13",
X"77",
X"13",
X"9d",
X"4a",
X"15",
X"c1",
X"a1",
X"41",
X"c3",
X"12",
X"fe",
X"01",
X"7d",
X"c1",
X"9e",
X"42",
X"cf",
X"20",
X"fd",
X"52",
X"21",
X"0f",
X"20",
X"6e",
X"44",
X"0c",
X"f1",
X"4c",
X"01",
X"aa",
X"35",
X"d9",
X"34",
X"ee",
X"20",
X"08",
X"b3",
X"37",
X"32",
X"43",
X"04",
X"4e",
X"21",
X"53",
X"20",
X"7c",
X"01",
X"97",
X"21",
X"b7",
X"07",
X"9c",
X"81",
X"e7",
X"42",
X"5f",
X"b3",
X"97",
X"63",
X"ac",
X"02",
X"c5",
X"41",
X"49",
X"e0",
X"58",
X"61",
X"76",
X"64",
X"85",
X"65",
X"94",
X"66",
X"a4",
X"22",
X"a6",
X"03",
X"c8",
X"22",
X"dc",
X"02",
X"68",
X"f2",
X"96",
X"42",
X"13",
X"82",
X"17",
X"02",
X"af",
X"34",
X"f6",
X"21",
X"fc",
X"06",
X"26",
X"80",
X"2a",
X"24",
X"36",
X"01",
X"8c",
X"00",
X"ff",
X"35",
X"4e",
X"a0",
X"55",
X"21",
X"77",
X"20",
X"87",
X"07",
X"89",
X"22",
X"ae",
X"21",
X"4c",
X"82",
X"9f",
X"34",
X"ec",
X"01",
X"03",
X"e7",
X"13",
X"67",
X"8d",
X"4a",
X"ad",
X"41",
X"0f",
X"a6",
X"fd",
X"10",
X"51",
X"4c",
X"00",
X"c7",
X"12",
X"c6",
X"42",
X"03",
X"92",
X"02",
X"42",
X"29",
X"12",
X"63",
X"12",
X"62",
X"42",
X"69",
X"14",
X"a5",
X"12",
X"a4",
X"42",
X"e2",
X"14",
X"e1",
X"44",
X"f8",
X"16",
X"37",
X"c1",
X"8f",
X"38",
X"02",
X"bb",
X"28",
X"7a",
X"68",
X"7a",
X"a8",
X"7a",
X"e0",
X"6a",
X"f0",
X"6a",
X"6d",
X"c5",
X"fd",
X"92",
X"31",
X"0f",
X"20",
X"6e",
X"40",
X"0d",
X"02",
X"37",
X"73",
X"ec",
X"00",
X"0c",
X"80",
X"3c",
X"00",
X"6c",
X"00",
X"9c",
X"00",
X"06",
X"c0",
X"c7",
X"73",
X"06",
X"83",
X"28",
X"72",
X"96",
X"40",
X"e7",
X"73",
X"26",
X"c0",
X"87",
X"7b",
X"d2",
X"41",
X"39",
X"f1",
X"c8",
X"f2",
X"97",
X"e3",
X"a3",
X"23",
X"e7",
X"02",
X"e3",
X"07",
X"f3",
X"22",
X"37",
X"e3",
X"9c",
X"00",
X"bc",
X"00",
X"ec",
X"00",
X"0c",
X"80",
X"3c",
X"00",
X"86",
X"21",
X"a6",
X"06",
X"b6",
X"24",
X"5c",
X"80",
X"7c",
X"00",
X"9c",
X"00",
X"29",
X"e1",
X"dc",
X"05",
X"f6",
X"41",
X"dc",
X"80",
X"e8",
X"72",
X"0c",
X"81",
X"27",
X"73",
X"4c",
X"01",
X"66",
X"74",
X"0d",
X"11",
X"3f",
X"35",
X"b6",
X"41",
X"2c",
X"82",
X"36",
X"40",
X"7c",
X"02",
X"86",
X"40",
X"f9",
X"61",
X"39",
X"e1",
X"ac",
X"04",
X"c6",
X"41",
X"0c",
X"83",
X"16",
X"41",
X"88",
X"f2",
X"39",
X"f1",
X"7c",
X"00",
X"89",
X"61",
X"9c",
X"00",
X"a7",
X"63",
X"bc",
X"00",
X"c5",
X"65",
X"dc",
X"00",
X"e3",
X"67",
X"f3",
X"67",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"55",
X"b1",
X"0f",
X"26",
X"cf",
X"33",
X"07",
X"b2",
X"15",
X"11",
X"52",
X"42",
X"99",
X"0b",
X"ac",
X"02",
X"d3",
X"24",
X"d6",
X"42",
X"d7",
X"25",
X"23",
X"84",
X"cf",
X"33",
X"07",
X"e3",
X"19",
X"61",
X"78",
X"7a",
X"ef",
X"33",
X"2c",
X"81",
X"46",
X"64",
X"55",
X"65",
X"65",
X"65",
X"ec",
X"74",
X"47",
X"82",
X"53",
X"05",
X"63",
X"21",
X"62",
X"41",
X"96",
X"22",
X"9a",
X"41",
X"cc",
X"03",
X"b9",
X"91",
X"39",
X"f1",
X"63",
X"26",
X"67",
X"27",
X"d3",
X"06",
X"fc",
X"01",
X"18",
X"e2",
X"d9",
X"07",
X"e9",
X"04",
X"0c",
X"86",
X"37",
X"22",
X"93",
X"24",
X"87",
X"84",
X"ac",
X"02",
X"c2",
X"41",
X"c3",
X"23",
X"d9",
X"71",
X"fc",
X"01",
X"7f",
X"b1",
X"9c",
X"00",
X"a7",
X"63",
X"b6",
X"64",
X"cc",
X"00",
X"d4",
X"66",
X"e3",
X"67",
X"f3",
X"67",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"50",
X"b1",
X"0f",
X"26",
X"fc",
X"00",
X"1f",
X"b3",
X"5c",
X"00",
X"65",
X"65",
X"74",
X"66",
X"83",
X"67",
X"93",
X"67",
X"dc",
X"73",
X"4c",
X"80",
X"b3",
X"20",
X"c9",
X"0b",
X"c3",
X"08",
X"d3",
X"2f",
X"dc",
X"00",
X"2c",
X"80",
X"4c",
X"00",
X"8c",
X"00",
X"d3",
X"2e",
X"ed",
X"4a",
X"fc",
X"00",
X"d7",
X"a1",
X"ec",
X"01",
X"4c",
X"80",
X"59",
X"11",
X"d8",
X"11",
X"da",
X"10",
X"37",
X"a0",
X"47",
X"04",
X"99",
X"11",
X"e7",
X"21",
X"3a",
X"90",
X"67",
X"20",
X"76",
X"10",
X"77",
X"60",
X"87",
X"07",
X"d8",
X"12",
X"39",
X"f1",
X"ac",
X"00",
X"e9",
X"71",
X"0c",
X"80",
X"2c",
X"00",
X"4c",
X"05",
X"c7",
X"7b",
X"39",
X"f1",
X"ec",
X"00",
X"f9",
X"11",
X"0c",
X"82",
X"6f",
X"34",
X"f8",
X"11",
X"fa",
X"10",
X"7f",
X"b2",
X"ac",
X"00",
X"b6",
X"64",
X"cc",
X"01",
X"e3",
X"67",
X"f3",
X"67",
X"8d",
X"c1",
X"cf",
X"26",
X"fd",
X"52",
X"b1",
X"0f",
X"20",
X"6e",
X"45",
X"39",
X"91",
X"b3",
X"04",
X"c3",
X"21",
X"c8",
X"11",
X"ca",
X"10",
X"49",
X"91",
X"7c",
X"73",
X"e8",
X"12",
X"88",
X"91",
X"8a",
X"10",
X"e7",
X"21",
X"05",
X"91",
X"07",
X"30",
X"17",
X"07",
X"27",
X"20",
X"49",
X"11",
X"9c",
X"01",
X"c8",
X"72",
X"23",
X"a6",
X"27",
X"26",
X"d3",
X"03",
X"d8",
X"7a",
X"89",
X"91",
X"d8",
X"72",
X"39",
X"f1",
X"a9",
X"11",
X"09",
X"f1",
X"63",
X"24",
X"67",
X"24",
X"d8",
X"62",
X"28",
X"91",
X"2a",
X"10",
X"56",
X"21",
X"70",
X"04",
X"79",
X"0b",
X"8c",
X"00",
X"94",
X"21",
X"9f",
X"35",
X"2f",
X"b8",
X"3d",
X"c1",
X"7f",
X"26",
X"fd",
X"06",
X"c1",
X"4c",
X"00",
X"f4",
X"4f",
X"0d",
X"02",
X"06",
X"20",
X"24",
X"4f",
X"35",
X"a0",
X"36",
X"20",
X"53",
X"46",
X"d5",
X"20",
X"d6",
X"20",
X"34",
X"a1",
X"73",
X"49",
X"74",
X"20",
X"94",
X"20",
X"b4",
X"20",
X"d4",
X"20",
X"f4",
X"20",
X"2e",
X"80",
X"59",
X"42",
X"4d",
X"c7",
X"fd",
X"96",
X"31",
X"0f",
X"26",
X"0d",
X"03",
X"1a",
X"60",
X"77",
X"42",
X"c4",
X"00",
X"c8",
X"62",
X"b9",
X"e1",
X"d3",
X"06",
X"d7",
X"07",
X"f9",
X"61",
X"0c",
X"81",
X"4e",
X"b1",
X"8e",
X"b1",
X"bc",
X"01",
X"e4",
X"50",
X"e9",
X"61",
X"0c",
X"81",
X"0d",
X"0a",
X"84",
X"43",
X"98",
X"72",
X"0d",
X"0c",
X"0f",
X"38",
X"1d",
X"c1",
X"5f",
X"26",
X"fd",
X"48",
X"0f",
X"0e",
X"01",
X"5e",
X"02",
X"a7",
X"00",
X"bc",
X"73",
X"1a",
X"e0",
X"39",
X"61",
X"58",
X"62",
X"77",
X"63",
X"97",
X"63",
X"b8",
X"62",
X"d6",
X"07",
X"f8",
X"62",
X"19",
X"e1",
X"75",
X"52",
X"86",
X"40",
X"87",
X"50",
X"95",
X"52",
X"93",
X"43",
X"a5",
X"21",
X"c5",
X"52",
X"d6",
X"40",
X"d7",
X"20",
X"e5",
X"06",
X"e6",
X"51",
X"3e",
X"8d",
X"5e",
X"03",
X"67",
X"52",
X"77",
X"52",
X"7e",
X"02",
X"9e",
X"03",
X"a6",
X"43",
X"a7",
X"23",
X"de",
X"05",
X"fe",
X"02",
X"1e",
X"83",
X"33",
X"54",
X"46",
X"40",
X"47",
X"21",
X"56",
X"04",
X"5e",
X"02",
X"83",
X"54",
X"93",
X"52",
X"96",
X"07",
X"97",
X"50",
X"be",
X"03",
X"c7",
X"23",
X"fe",
X"02",
X"0c",
X"82",
X"43",
X"45",
X"45",
X"24",
X"46",
X"24",
X"90",
X"08",
X"95",
X"51",
X"78",
X"fa",
X"d7",
X"73",
X"39",
X"f1",
X"8c",
X"01",
X"a8",
X"52",
X"b8",
X"52",
X"cc",
X"01",
X"5f",
X"b3",
X"97",
X"63",
X"9e",
X"00",
X"0e",
X"81",
X"16",
X"24",
X"66",
X"04",
X"8e",
X"00",
X"fe",
X"01",
X"08",
X"d2",
X"0e",
X"06",
X"6f",
X"47",
X"9e",
X"0f",
X"0e",
X"82",
X"2d",
X"47",
X"28",
X"7a",
X"68",
X"7a",
X"a8",
X"7a",
X"ae",
X"01",
X"de",
X"0f",
X"6d",
X"c5",
X"fd",
X"48",
X"0f",
X"0e",
X"01",
X"5e",
X"02",
X"bc",
X"01",
X"fc",
X"01",
X"2c",
X"82",
X"41",
X"52",
X"4e",
X"04",
X"67",
X"25",
X"68",
X"24",
X"69",
X"24",
X"ba",
X"42",
X"c7",
X"04",
X"de",
X"0b",
X"b2",
X"87",
X"fe",
X"02",
X"2c",
X"e1",
X"2c",
X"71",
X"67",
X"01",
X"77",
X"00",
X"87",
X"01",
X"8e",
X"00",
X"ee",
X"01",
X"f6",
X"02",
X"03",
X"85",
X"05",
X"02",
X"13",
X"21",
X"16",
X"02",
X"27",
X"02",
X"2e",
X"02",
X"88",
X"72",
X"c7",
X"20",
X"d7",
X"07",
X"e4",
X"76",
X"07",
X"a0",
X"17",
X"06",
X"48",
X"7a",
X"76",
X"20",
X"98",
X"72",
X"79",
X"e1",
X"88",
X"62",
X"9c",
X"01",
X"b7",
X"73",
X"dc",
X"01",
X"f8",
X"62",
X"fe",
X"01",
X"08",
X"e2",
X"0e",
X"00",
X"6e",
X"02",
X"73",
X"20",
X"77",
X"23",
X"83",
X"04",
X"93",
X"20",
X"ae",
X"00",
X"fe",
X"0a",
X"0e",
X"82",
X"39",
X"71",
X"a8",
X"72",
X"e7",
X"73",
X"0c",
X"81",
X"8f",
X"32",
X"ae",
X"00",
X"fe",
X"04",
X"04",
X"d1",
X"17",
X"04",
X"26",
X"49",
X"27",
X"29",
X"df",
X"33",
X"fe",
X"02",
X"44",
X"f6",
X"7c",
X"01",
X"8e",
X"06",
X"bf",
X"47",
X"ee",
X"0f",
X"4d",
X"c7",
X"0e",
X"82",
X"68",
X"7a",
X"ae",
X"01",
X"de",
X"0f",
X"6d",
X"c5",
X"fd",
X"48",
X"01",
X"0e",
X"01",
X"00",
X"5a",
X"3e",
X"06",
X"45",
X"46",
X"47",
X"46",
X"53",
X"44",
X"ae",
X"01",
X"df",
X"4a",
X"4d",
X"c7",
X"0e",
X"81",
X"00",
X"5a",
X"2e",
X"04",
X"37",
X"28",
X"3a",
X"48",
X"46",
X"47",
X"c7",
X"07",
X"ce",
X"0f",
X"df",
X"4a",
X"4d",
X"c7",
X"0e",
X"81",
X"00",
X"5a",
X"33",
X"53",
X"43",
X"51",
X"46",
X"40",
X"47",
X"50",
X"53",
X"04",
X"55",
X"40",
X"56",
X"50",
X"62",
X"43",
X"64",
X"40",
X"65",
X"50",
X"71",
X"41",
X"73",
X"51",
X"83",
X"51",
X"94",
X"40",
X"95",
X"50",
X"a3",
X"50",
X"a5",
X"40",
X"a6",
X"50",
X"b3",
X"51",
X"b6",
X"40",
X"b7",
X"50",
X"c3",
X"53",
X"df",
X"4a",
X"4d",
X"c7",
X"0e",
X"81",
X"00",
X"5a",
X"2e",
X"02",
X"36",
X"47",
X"37",
X"52",
X"3a",
X"49",
X"47",
X"25",
X"a7",
X"52",
X"d7",
X"04",
X"df",
X"4a",
X"4d",
X"c7",
X"0e",
X"81",
X"00",
X"5a",
X"3e",
X"02",
X"44",
X"51",
X"53",
X"44",
X"54",
X"44",
X"55",
X"24",
X"a1",
X"54",
X"ae",
X"01",
X"b4",
X"21",
X"df",
X"4a",
X"e5",
X"07",
X"4d",
X"c7",
X"fd",
X"41",
X"01",
X"b4",
X"34",
X"c8",
X"52",
X"f2",
X"51",
X"47",
X"d3",
X"6c",
X"03",
X"65",
X"49",
X"9e",
X"07",
X"be",
X"01",
X"cc",
X"03",
X"fe",
X"07",
X"0d",
X"c9",
X"1e",
X"01",
X"6c",
X"01",
X"62",
X"35",
X"63",
X"53",
X"8a",
X"41",
X"ac",
X"01",
X"b3",
X"53",
X"e9",
X"51",
X"26",
X"c3",
X"27",
X"33",
X"63",
X"43",
X"64",
X"33",
X"ba",
X"60",
X"c9",
X"61",
X"ce",
X"0b",
X"e5",
X"09",
X"ee",
X"0f",
X"7d",
X"ca",
X"7d",
X"47",
X"fd",
X"41",
X"01",
X"b8",
X"52",
X"ea",
X"41",
X"27",
X"b2",
X"b3",
X"42",
X"16",
X"d4",
X"4a",
X"42",
X"a5",
X"51",
X"a7",
X"31",
X"27",
X"d3",
X"08",
X"e2",
X"16",
X"64",
X"2c",
X"04",
X"38",
X"42",
X"76",
X"64",
X"88",
X"62",
X"de",
X"07",
X"fe",
X"01",
X"0d",
X"c9",
X"23",
X"32",
X"31",
X"51",
X"98",
X"52",
X"0d",
X"c9",
X"59",
X"42",
X"63",
X"53",
X"67",
X"31",
X"14",
X"c2",
X"36",
X"31",
X"87",
X"53",
X"17",
X"e3",
X"29",
X"61",
X"30",
X"62",
X"3c",
X"08",
X"42",
X"37",
X"59",
X"40",
X"6a",
X"42",
X"99",
X"40",
X"c9",
X"61",
X"d7",
X"63",
X"39",
X"d1",
X"58",
X"52",
X"c3",
X"67",
X"d3",
X"31",
X"dc",
X"06",
X"f7",
X"42",
X"fa",
X"42",
X"23",
X"b1",
X"43",
X"67",
X"c3",
X"34",
X"c7",
X"34",
X"d1",
X"51",
X"43",
X"b3",
X"47",
X"33",
X"9a",
X"30",
X"a9",
X"61",
X"b8",
X"62",
X"be",
X"0b",
X"d5",
X"09",
X"de",
X"0f",
X"0d",
X"ca",
X"7d",
X"47",
X"fd",
X"49",
X"0f",
X"1e",
X"01",
X"39",
X"73",
X"5e",
X"07",
X"ae",
X"0b",
X"1e",
X"82",
X"6e",
X"88",
X"9e",
X"02",
X"0d",
X"04",
X"2e",
X"0b",
X"45",
X"09",
X"4e",
X"0f",
X"ed",
X"47",
X"fd",
X"ff",
X"ad",
X"72",
X"07",
X"20",
X"04",
X"8e",
X"e4",
X"8f",
X"67",
X"85",
X"71",
X"90",
X"ea",
X"ae",
X"ae",
X"53",
X"07",
X"bd",
X"fc",
X"06",
X"8d",
X"fc",
X"06",
X"20",
X"4a",
X"b0",
X"ad",
X"72",
X"07",
X"c9",
X"03",
X"b0",
X"01",
X"60",
X"20",
X"24",
X"b6",
X"a2",
X"00",
X"86",
X"08",
X"20",
X"47",
X"c0",
X"20",
X"c3",
X"84",
X"e8",
X"e0",
X"06",
X"d0",
X"f3",
X"20",
X"80",
X"f1",
X"20",
X"2a",
X"f1",
X"20",
X"e9",
X"ee",
X"20",
X"d4",
X"be",
X"a2",
X"01",
X"86",
X"08",
X"20",
X"70",
X"be",
X"ca",
X"86",
X"08",
X"20",
X"70",
X"be",
X"20",
X"96",
X"bb",
X"20",
X"bc",
X"b9",
X"20",
X"b8",
X"b7",
X"20",
X"55",
X"b8",
X"20",
X"4f",
X"b7",
X"20",
X"e1",
X"89",
X"a5",
X"b5",
X"c9",
X"02",
X"10",
X"11",
X"ad",
X"9f",
X"07",
X"f0",
X"1e",
X"c9",
X"04",
X"d0",
X"08",
X"ad",
X"7f",
X"07",
X"d0",
X"03",
X"20",
X"ed",
X"90",
X"ac",
X"9f",
X"07",
X"a5",
X"09",
X"c0",
X"08",
X"b0",
X"02",
X"4a",
X"4a",
X"4a",
X"20",
X"88",
X"b2",
X"4c",
X"67",
X"af",
X"20",
X"9a",
X"b2",
X"a5",
X"0a",
X"85",
X"0d",
X"a9",
X"00",
X"85",
X"0c",
X"ad",
X"73",
X"07",
X"c9",
X"06",
X"f0",
X"1c",
X"ad",
X"1f",
X"07",
X"d0",
X"14",
X"ad",
X"3d",
X"07",
X"c9",
X"20",
X"30",
X"10",
X"ad",
X"3d",
X"07",
X"e9",
X"20",
X"8d",
X"3d",
X"07",
X"a9",
X"00",
X"8d",
X"40",
X"03",
X"20",
X"b0",
X"92",
X"60",
X"ad",
X"ff",
X"06",
X"18",
X"6d",
X"a1",
X"03",
X"8d",
X"ff",
X"06",
X"ad",
X"23",
X"07",
X"d0",
X"59",
X"ad",
X"55",
X"07",
X"c9",
X"50",
X"90",
X"52",
X"ad",
X"85",
X"07",
X"d0",
X"4d",
X"ac",
X"ff",
X"06",
X"88",
X"30",
X"47",
X"c8",
X"c0",
X"02",
X"90",
X"01",
X"88",
X"ad",
X"55",
X"07",
X"c9",
X"70",
X"90",
X"03",
X"ac",
X"ff",
X"06",
X"98",
X"8d",
X"75",
X"07",
X"18",
X"6d",
X"3d",
X"07",
X"8d",
X"3d",
X"07",
X"98",
X"18",
X"6d",
X"1c",
X"07",
X"8d",
X"1c",
X"07",
X"8d",
X"3f",
X"07",
X"ad",
X"1a",
X"07",
X"69",
X"00",
X"8d",
X"1a",
X"07",
X"29",
X"01",
X"85",
X"00",
X"ad",
X"78",
X"07",
X"29",
X"fe",
X"05",
X"00",
X"8d",
X"78",
X"07",
X"20",
X"38",
X"b0",
X"a9",
X"08",
X"8d",
X"95",
X"07",
X"4c",
X"00",
X"b0",
X"a9",
X"00",
X"8d",
X"75",
X"07",
X"a2",
X"00",
X"20",
X"f6",
X"f1",
X"85",
X"00",
X"a0",
X"00",
X"0a",
X"b0",
X"07",
X"c8",
X"a5",
X"00",
X"29",
X"20",
X"f0",
X"1b",
X"b9",
X"1c",
X"07",
X"38",
X"f9",
X"34",
X"b0",
X"85",
X"86",
X"b9",
X"1a",
X"07",
X"e9",
X"00",
X"85",
X"6d",
X"a5",
X"0c",
X"d9",
X"36",
X"b0",
X"f0",
X"04",
X"a9",
X"00",
X"85",
X"57",
X"a9",
X"00",
X"8d",
X"a1",
X"03",
X"60",
X"00",
X"10",
X"01",
X"02",
X"ad",
X"1c",
X"07",
X"18",
X"69",
X"ff",
X"8d",
X"1d",
X"07",
X"ad",
X"1a",
X"07",
X"69",
X"00",
X"8d",
X"1b",
X"07",
X"60",
X"a5",
X"0e",
X"20",
X"04",
X"8e",
X"31",
X"91",
X"c7",
X"b1",
X"06",
X"b2",
X"e5",
X"b1",
X"a4",
X"b2",
X"ca",
X"b2",
X"cd",
X"91",
X"69",
X"b0",
X"e9",
X"b0",
X"33",
X"b2",
X"45",
X"b2",
X"69",
X"b2",
X"7d",
X"b2",
X"ad",
X"52",
X"07",
X"c9",
X"02",
X"f0",
X"2b",
X"a9",
X"00",
X"a4",
X"ce",
X"c0",
X"30",
X"90",
X"6e",
X"ad",
X"10",
X"07",
X"c9",
X"06",
X"f0",
X"04",
X"c9",
X"07",
X"d0",
X"50",
X"ad",
X"c4",
X"03",
X"d0",
X"05",
X"a9",
X"01",
X"4c",
X"e6",
X"b0",
X"20",
X"1f",
X"b2",
X"ce",
X"de",
X"06",
X"d0",
X"50",
X"ee",
X"69",
X"07",
X"4c",
X"15",
X"b3",
X"ad",
X"58",
X"07",
X"d0",
X"0c",
X"a9",
X"ff",
X"20",
X"00",
X"b2",
X"a5",
X"ce",
X"c9",
X"91",
X"90",
X"28",
X"60",
X"ad",
X"99",
X"03",
X"c9",
X"60",
X"d0",
X"32",
X"a5",
X"ce",
X"c9",
X"99",
X"a0",
X"00",
X"a9",
X"01",
X"90",
X"0a",
X"a9",
X"03",
X"85",
X"1d",
X"c8",
X"a9",
X"08",
X"8d",
X"b4",
X"05",
X"8c",
X"16",
X"07",
X"20",
X"e6",
X"b0",
X"a5",
X"86",
X"c9",
X"48",
X"90",
X"12",
X"a9",
X"08",
X"85",
X"0e",
X"a9",
X"01",
X"85",
X"33",
X"4a",
X"8d",
X"52",
X"07",
X"8d",
X"16",
X"07",
X"8d",
X"58",
X"07",
X"60",
X"8d",
X"fc",
X"06",
X"a5",
X"0e",
X"c9",
X"0b",
X"f0",
X"3c",
X"ad",
X"4e",
X"07",
X"d0",
X"10",
X"a4",
X"b5",
X"88",
X"d0",
X"06",
X"a5",
X"ce",
X"c9",
X"d0",
X"90",
X"05",
X"a9",
X"00",
X"8d",
X"fc",
X"06",
X"ad",
X"fc",
X"06",
X"29",
X"c0",
X"85",
X"0a",
X"ad",
X"fc",
X"06",
X"29",
X"03",
X"85",
X"0c",
X"ad",
X"fc",
X"06",
X"29",
X"0c",
X"85",
X"0b",
X"29",
X"04",
X"f0",
X"0e",
X"a5",
X"1d",
X"d0",
X"0a",
X"a4",
X"0c",
X"f0",
X"06",
X"a9",
X"00",
X"85",
X"0c",
X"85",
X"0b",
X"20",
X"29",
X"b3",
X"a0",
X"01",
X"ad",
X"54",
X"07",
X"d0",
X"09",
X"a0",
X"00",
X"ad",
X"14",
X"07",
X"f0",
X"02",
X"a0",
X"02",
X"8c",
X"99",
X"04",
X"a9",
X"01",
X"a4",
X"57",
X"f0",
X"05",
X"10",
X"01",
X"0a",
X"85",
X"45",
X"20",
X"93",
X"af",
X"20",
X"80",
X"f1",
X"20",
X"2a",
X"f1",
X"a2",
X"00",
X"20",
X"9c",
X"e2",
X"20",
X"64",
X"dc",
X"a5",
X"ce",
X"c9",
X"40",
X"90",
X"16",
X"a5",
X"0e",
X"c9",
X"05",
X"f0",
X"10",
X"c9",
X"07",
X"f0",
X"0c",
X"c9",
X"04",
X"90",
X"08",
X"ad",
X"c4",
X"03",
X"29",
X"df",
X"8d",
X"c4",
X"03",
X"a5",
X"b5",
X"c9",
X"02",
X"30",
X"3b",
X"a2",
X"01",
X"8e",
X"23",
X"07",
X"a0",
X"04",
X"84",
X"07",
X"a2",
X"00",
X"ac",
X"59",
X"07",
X"d0",
X"05",
X"ac",
X"43",
X"07",
X"d0",
X"16",
X"e8",
X"a4",
X"0e",
X"c0",
X"0b",
X"f0",
X"0f",
X"ac",
X"12",
X"07",
X"d0",
X"06",
X"c8",
X"84",
X"fc",
X"8c",
X"12",
X"07",
X"a0",
X"06",
X"84",
X"07",
X"c5",
X"07",
X"30",
X"0c",
X"ca",
X"30",
X"0a",
X"ac",
X"b1",
X"07",
X"d0",
X"04",
X"a9",
X"06",
X"85",
X"0e",
X"60",
X"a9",
X"00",
X"8d",
X"58",
X"07",
X"20",
X"dd",
X"b1",
X"ee",
X"52",
X"07",
X"60",
X"a5",
X"b5",
X"d0",
X"06",
X"a5",
X"ce",
X"c9",
X"e4",
X"90",
X"0c",
X"a9",
X"08",
X"8d",
X"58",
X"07",
X"a0",
X"03",
X"84",
X"1d",
X"4c",
X"e6",
X"b0",
X"a9",
X"02",
X"8d",
X"52",
X"07",
X"4c",
X"13",
X"b2",
X"a9",
X"01",
X"20",
X"00",
X"b2",
X"20",
X"93",
X"af",
X"a0",
X"00",
X"ad",
X"d6",
X"06",
X"d0",
X"17",
X"c8",
X"ad",
X"4e",
X"07",
X"c9",
X"03",
X"d0",
X"0f",
X"c8",
X"4c",
X"0b",
X"b2",
X"18",
X"65",
X"ce",
X"85",
X"ce",
X"60",
X"20",
X"1f",
X"b2",
X"a0",
X"02",
X"ce",
X"de",
X"06",
X"d0",
X"0e",
X"8c",
X"52",
X"07",
X"ee",
X"74",
X"07",
X"a9",
X"00",
X"8d",
X"72",
X"07",
X"8d",
X"22",
X"07",
X"60",
X"a9",
X"08",
X"85",
X"57",
X"a0",
X"01",
X"a5",
X"86",
X"29",
X"0f",
X"d0",
X"03",
X"85",
X"57",
X"a8",
X"98",
X"20",
X"e6",
X"b0",
X"60",
X"ad",
X"47",
X"07",
X"c9",
X"f8",
X"d0",
X"03",
X"4c",
X"55",
X"b2",
X"c9",
X"c4",
X"d0",
X"03",
X"20",
X"73",
X"b2",
X"60",
X"ad",
X"47",
X"07",
X"c9",
X"f0",
X"b0",
X"07",
X"c9",
X"c8",
X"f0",
X"23",
X"4c",
X"e9",
X"b0",
X"d0",
X"13",
X"ac",
X"0b",
X"07",
X"d0",
X"0e",
X"8c",
X"0d",
X"07",
X"ee",
X"0b",
X"07",
X"ad",
X"54",
X"07",
X"49",
X"01",
X"8d",
X"54",
X"07",
X"60",
X"ad",
X"47",
X"07",
X"c9",
X"f0",
X"b0",
X"33",
X"4c",
X"e9",
X"b0",
X"a9",
X"00",
X"8d",
X"47",
X"07",
X"a9",
X"08",
X"85",
X"0e",
X"60",
X"ad",
X"47",
X"07",
X"c9",
X"c0",
X"f0",
X"13",
X"a5",
X"09",
X"4a",
X"4a",
X"29",
X"03",
X"85",
X"00",
X"ad",
X"c4",
X"03",
X"29",
X"fc",
X"05",
X"00",
X"8d",
X"c4",
X"03",
X"60",
X"20",
X"73",
X"b2",
X"ad",
X"c4",
X"03",
X"29",
X"fc",
X"8d",
X"c4",
X"03",
X"60",
X"60",
X"a5",
X"1b",
X"c9",
X"30",
X"d0",
X"15",
X"ad",
X"13",
X"07",
X"85",
X"ff",
X"a9",
X"00",
X"8d",
X"13",
X"07",
X"a4",
X"ce",
X"c0",
X"9e",
X"b0",
X"02",
X"a9",
X"04",
X"4c",
X"e6",
X"b0",
X"e6",
X"0e",
X"60",
X"15",
X"23",
X"16",
X"1b",
X"17",
X"18",
X"23",
X"63",
X"a9",
X"01",
X"20",
X"e6",
X"b0",
X"a5",
X"ce",
X"c9",
X"ae",
X"90",
X"0e",
X"ad",
X"23",
X"07",
X"f0",
X"09",
X"a9",
X"20",
X"85",
X"fc",
X"a9",
X"00",
X"8d",
X"23",
X"07",
X"ad",
X"90",
X"04",
X"4a",
X"b0",
X"0d",
X"ad",
X"46",
X"07",
X"d0",
X"03",
X"ee",
X"46",
X"07",
X"a9",
X"20",
X"8d",
X"c4",
X"03",
X"ad",
X"46",
X"07",
X"c9",
X"05",
X"d0",
X"2b",
X"ee",
X"5c",
X"07",
X"ad",
X"5c",
X"07",
X"c9",
X"03",
X"d0",
X"0e",
X"ac",
X"5f",
X"07",
X"ad",
X"48",
X"07",
X"d9",
X"c2",
X"b2",
X"90",
X"03",
X"ee",
X"5d",
X"07",
X"ee",
X"60",
X"07",
X"20",
X"03",
X"9c",
X"ee",
X"57",
X"07",
X"20",
X"13",
X"b2",
X"8d",
X"5b",
X"07",
X"a9",
X"80",
X"85",
X"fc",
X"60",
X"a9",
X"00",
X"ac",
X"54",
X"07",
X"d0",
X"08",
X"a5",
X"1d",
X"d0",
X"07",
X"a5",
X"0b",
X"29",
X"04",
X"8d",
X"14",
X"07",
X"20",
X"50",
X"b4",
X"ad",
X"0b",
X"07",
X"d0",
X"16",
X"a5",
X"1d",
X"c9",
X"03",
X"f0",
X"05",
X"a0",
X"18",
X"8c",
X"89",
X"07",
X"20",
X"04",
X"8e",
X"5a",
X"b3",
X"76",
X"b3",
X"6d",
X"b3",
X"cf",
X"b3",
X"60",
X"20",
X"8f",
X"b5",
X"a5",
X"0c",
X"f0",
X"02",
X"85",
X"33",
X"20",
X"cc",
X"b5",
X"20",
X"09",
X"bf",
X"8d",
X"ff",
X"06",
X"60",
X"ad",
X"0a",
X"07",
X"8d",
X"09",
X"07",
X"4c",
X"ac",
X"b3",
X"a4",
X"9f",
X"10",
X"13",
X"a5",
X"0a",
X"29",
X"80",
X"25",
X"0d",
X"d0",
X"11",
X"ad",
X"08",
X"07",
X"38",
X"e5",
X"ce",
X"cd",
X"06",
X"07",
X"90",
X"06",
X"ad",
X"0a",
X"07",
X"8d",
X"09",
X"07",
X"ad",
X"04",
X"07",
X"f0",
X"14",
X"20",
X"8f",
X"b5",
X"a5",
X"ce",
X"c9",
X"14",
X"b0",
X"05",
X"a9",
X"18",
X"8d",
X"09",
X"07",
X"a5",
X"0c",
X"f0",
X"02",
X"85",
X"33",
X"a5",
X"0c",
X"f0",
X"03",
X"20",
X"cc",
X"b5",
X"20",
X"09",
X"bf",
X"8d",
X"ff",
X"06",
X"a5",
X"0e",
X"c9",
X"0b",
X"d0",
X"05",
X"a9",
X"28",
X"8d",
X"09",
X"07",
X"4c",
X"4d",
X"bf",
X"0e",
X"04",
X"fc",
X"f2",
X"00",
X"00",
X"ff",
X"ff",
X"ad",
X"16",
X"04",
X"18",
X"6d",
X"33",
X"04",
X"8d",
X"16",
X"04",
X"a0",
X"00",
X"a5",
X"9f",
X"10",
X"01",
X"88",
X"84",
X"00",
X"65",
X"ce",
X"85",
X"ce",
X"a5",
X"b5",
X"65",
X"00",
X"85",
X"b5",
X"a5",
X"0c",
X"2d",
X"90",
X"04",
X"f0",
X"2d",
X"ac",
X"89",
X"07",
X"d0",
X"27",
X"a0",
X"18",
X"8c",
X"89",
X"07",
X"a2",
X"00",
X"a4",
X"33",
X"4a",
X"b0",
X"02",
X"e8",
X"e8",
X"88",
X"f0",
X"01",
X"e8",
X"a5",
X"86",
X"18",
X"7d",
X"c7",
X"b3",
X"85",
X"86",
X"a5",
X"6d",
X"7d",
X"cb",
X"b3",
X"85",
X"6d",
X"a5",
X"0c",
X"49",
X"03",
X"85",
X"33",
X"60",
X"8d",
X"89",
X"07",
X"60",
X"20",
X"20",
X"1e",
X"28",
X"28",
X"0d",
X"04",
X"70",
X"70",
X"60",
X"90",
X"90",
X"0a",
X"09",
X"fc",
X"fc",
X"fc",
X"fb",
X"fb",
X"fe",
X"ff",
X"00",
X"00",
X"00",
X"00",
X"00",
X"80",
X"00",
X"d8",
X"e8",
X"f0",
X"28",
X"18",
X"10",
X"0c",
X"e4",
X"98",
X"d0",
X"00",
X"ff",
X"01",
X"00",
X"20",
X"ff",
X"a5",
X"1d",
X"c9",
X"03",
X"d0",
X"23",
X"a0",
X"00",
X"a5",
X"0b",
X"2d",
X"90",
X"04",
X"f0",
X"06",
X"c8",
X"29",
X"08",
X"d0",
X"01",
X"c8",
X"be",
X"4d",
X"b4",
X"8e",
X"33",
X"04",
X"a9",
X"08",
X"be",
X"4a",
X"b4",
X"86",
X"9f",
X"30",
X"01",
X"4a",
X"8d",
X"0c",
X"07",
X"60",
X"ad",
X"0e",
X"07",
X"d0",
X"0a",
X"a5",
X"0a",
X"29",
X"80",
X"f0",
X"04",
X"25",
X"0d",
X"f0",
X"03",
X"4c",
X"1c",
X"b5",
X"a5",
X"1d",
X"f0",
X"11",
X"ad",
X"04",
X"07",
X"f0",
X"f4",
X"ad",
X"82",
X"07",
X"d0",
X"07",
X"a5",
X"9f",
X"10",
X"03",
X"4c",
X"1c",
X"b5",
X"a9",
X"20",
X"8d",
X"82",
X"07",
X"a0",
X"00",
X"8c",
X"16",
X"04",
X"8c",
X"33",
X"04",
X"a5",
X"b5",
X"8d",
X"07",
X"07",
X"a5",
X"ce",
X"8d",
X"08",
X"07",
X"a9",
X"01",
X"85",
X"1d",
X"ad",
X"00",
X"07",
X"c9",
X"09",
X"90",
X"10",
X"c8",
X"c9",
X"10",
X"90",
X"0b",
X"c8",
X"c9",
X"19",
X"90",
X"06",
X"c8",
X"c9",
X"1c",
X"90",
X"01",
X"c8",
X"a9",
X"01",
X"8d",
X"06",
X"07",
X"ad",
X"04",
X"07",
X"f0",
X"08",
X"a0",
X"05",
X"ad",
X"7d",
X"04",
X"f0",
X"01",
X"c8",
X"b9",
X"24",
X"b4",
X"8d",
X"09",
X"07",
X"b9",
X"2b",
X"b4",
X"8d",
X"0a",
X"07",
X"b9",
X"39",
X"b4",
X"8d",
X"33",
X"04",
X"b9",
X"32",
X"b4",
X"85",
X"9f",
X"ad",
X"04",
X"07",
X"f0",
X"11",
X"a9",
X"04",
X"85",
X"ff",
X"a5",
X"ce",
X"c9",
X"14",
X"b0",
X"12",
X"a9",
X"00",
X"85",
X"9f",
X"4c",
X"1c",
X"b5",
X"a9",
X"01",
X"ac",
X"54",
X"07",
X"f0",
X"02",
X"a9",
X"80",
X"85",
X"ff",
X"a0",
X"00",
X"84",
X"00",
X"a5",
X"1d",
X"f0",
X"09",
X"ad",
X"00",
X"07",
X"c9",
X"19",
X"b0",
X"33",
X"90",
X"18",
X"c8",
X"ad",
X"4e",
X"07",
X"f0",
X"12",
X"88",
X"a5",
X"0c",
X"c5",
X"45",
X"d0",
X"0b",
X"a5",
X"0a",
X"29",
X"40",
X"d0",
X"19",
X"ad",
X"83",
X"07",
X"d0",
X"19",
X"c8",
X"e6",
X"00",
X"ad",
X"03",
X"07",
X"d0",
X"07",
X"ad",
X"00",
X"07",
X"c9",
X"21",
X"90",
X"0a",
X"e6",
X"00",
X"4c",
X"5e",
X"b5",
X"a9",
X"0a",
X"8d",
X"83",
X"07",
X"b9",
X"40",
X"b4",
X"8d",
X"50",
X"04",
X"a5",
X"0e",
X"c9",
X"07",
X"d0",
X"02",
X"a0",
X"03",
X"b9",
X"43",
X"b4",
X"8d",
X"56",
X"04",
X"a4",
X"00",
X"b9",
X"47",
X"b4",
X"8d",
X"02",
X"07",
X"a9",
X"00",
X"8d",
X"01",
X"07",
X"a5",
X"33",
X"c5",
X"45",
X"f0",
X"06",
X"0e",
X"02",
X"07",
X"2e",
X"01",
X"07",
X"60",
X"02",
X"04",
X"07",
X"a0",
X"00",
X"ad",
X"00",
X"07",
X"c9",
X"1c",
X"b0",
X"15",
X"c8",
X"c9",
X"0e",
X"b0",
X"01",
X"c8",
X"ad",
X"fc",
X"06",
X"29",
X"7f",
X"f0",
X"20",
X"29",
X"03",
X"c5",
X"45",
X"d0",
X"08",
X"a9",
X"00",
X"8d",
X"03",
X"07",
X"4c",
X"c5",
X"b5",
X"ad",
X"00",
X"07",
X"c9",
X"0b",
X"b0",
X"0b",
X"a5",
X"33",
X"85",
X"45",
X"a9",
X"00",
X"85",
X"57",
X"8d",
X"05",
X"07",
X"b9",
X"8c",
X"b5",
X"8d",
X"0c",
X"07",
X"60",
X"2d",
X"90",
X"04",
X"c9",
X"00",
X"d0",
X"08",
X"a5",
X"57",
X"f0",
X"49",
X"10",
X"23",
X"30",
X"03",
X"4a",
X"90",
X"1e",
X"ad",
X"05",
X"07",
X"18",
X"6d",
X"02",
X"07",
X"8d",
X"05",
X"07",
X"a5",
X"57",
X"6d",
X"01",
X"07",
X"85",
X"57",
X"cd",
X"56",
X"04",
X"30",
X"23",
X"ad",
X"56",
X"04",
X"85",
X"57",
X"4c",
X"20",
X"b6",
X"ad",
X"05",
X"07",
X"38",
X"ed",
X"02",
X"07",
X"8d",
X"05",
X"07",
X"a5",
X"57",
X"ed",
X"01",
X"07",
X"85",
X"57",
X"cd",
X"50",
X"04",
X"10",
X"05",
X"ad",
X"50",
X"04",
X"85",
X"57",
X"c9",
X"00",
X"10",
X"05",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"8d",
X"00",
X"07",
X"60",
X"ad",
X"56",
X"07",
X"c9",
X"02",
X"90",
X"43",
X"a5",
X"0a",
X"29",
X"40",
X"f0",
X"33",
X"25",
X"0d",
X"d0",
X"2f",
X"ad",
X"ce",
X"06",
X"29",
X"01",
X"aa",
X"b5",
X"24",
X"d0",
X"25",
X"a4",
X"b5",
X"88",
X"d0",
X"20",
X"ad",
X"14",
X"07",
X"d0",
X"1b",
X"a5",
X"1d",
X"c9",
X"03",
X"f0",
X"15",
X"a9",
X"20",
X"85",
X"ff",
X"a9",
X"02",
X"95",
X"24",
X"ac",
X"0c",
X"07",
X"8c",
X"11",
X"07",
X"88",
X"8c",
X"81",
X"07",
X"ee",
X"ce",
X"06",
X"a2",
X"00",
X"20",
X"89",
X"b6",
X"a2",
X"01",
X"20",
X"89",
X"b6",
X"ad",
X"4e",
X"07",
X"d0",
X"13",
X"a2",
X"02",
X"86",
X"08",
X"20",
X"f9",
X"b6",
X"20",
X"31",
X"f1",
X"20",
X"91",
X"f1",
X"20",
X"e1",
X"ed",
X"ca",
X"10",
X"ef",
X"60",
X"40",
X"c0",
X"86",
X"08",
X"b5",
X"24",
X"0a",
X"b0",
X"63",
X"b4",
X"24",
X"f0",
X"5e",
X"88",
X"f0",
X"27",
X"a5",
X"86",
X"69",
X"04",
X"95",
X"8d",
X"a5",
X"6d",
X"69",
X"00",
X"95",
X"74",
X"a5",
X"ce",
X"95",
X"d5",
X"a9",
X"01",
X"95",
X"bc",
X"a4",
X"33",
X"88",
X"b9",
X"87",
X"b6",
X"95",
X"5e",
X"a9",
X"04",
X"95",
X"a6",
X"a9",
X"07",
X"9d",
X"a0",
X"04",
X"d6",
X"24",
X"8a",
X"18",
X"69",
X"07",
X"aa",
X"a9",
X"50",
X"85",
X"00",
X"a9",
X"03",
X"85",
X"02",
X"a9",
X"00",
X"20",
X"d7",
X"bf",
X"20",
X"0f",
X"bf",
X"a6",
X"08",
X"20",
X"3b",
X"f1",
X"20",
X"87",
X"f1",
X"20",
X"2d",
X"e2",
X"20",
X"c8",
X"e1",
X"ad",
X"d2",
X"03",
X"29",
X"cc",
X"d0",
X"06",
X"20",
X"d9",
X"d6",
X"4c",
X"de",
X"ec",
X"a9",
X"00",
X"95",
X"24",
X"60",
X"20",
X"3b",
X"f1",
X"4c",
X"09",
X"ed",
X"bd",
X"a8",
X"07",
X"29",
X"01",
X"85",
X"07",
X"b5",
X"e4",
X"c9",
X"f8",
X"d0",
X"2c",
X"ad",
X"92",
X"07",
X"d0",
X"3f",
X"a0",
X"00",
X"a5",
X"33",
X"4a",
X"90",
X"02",
X"a0",
X"08",
X"98",
X"65",
X"86",
X"95",
X"9c",
X"a5",
X"6d",
X"69",
X"00",
X"95",
X"83",
X"a5",
X"ce",
X"18",
X"69",
X"08",
X"95",
X"e4",
X"a9",
X"01",
X"95",
X"cb",
X"a4",
X"07",
X"b9",
X"4d",
X"b7",
X"8d",
X"92",
X"07",
X"a4",
X"07",
X"bd",
X"2c",
X"04",
X"38",
X"f9",
X"4b",
X"b7",
X"9d",
X"2c",
X"04",
X"b5",
X"e4",
X"e9",
X"00",
X"c9",
X"20",
X"b0",
X"02",
X"a9",
X"f8",
X"95",
X"e4",
X"60",
X"ff",
X"50",
X"40",
X"20",
X"ad",
X"70",
X"07",
X"f0",
X"4f",
X"a5",
X"0e",
X"c9",
X"08",
X"90",
X"49",
X"c9",
X"0b",
X"f0",
X"45",
X"a5",
X"b5",
X"c9",
X"02",
X"b0",
X"3f",
X"ad",
X"87",
X"07",
X"d0",
X"3a",
X"ad",
X"f8",
X"07",
X"0d",
X"f9",
X"07",
X"0d",
X"fa",
X"07",
X"f0",
X"26",
X"ac",
X"f8",
X"07",
X"88",
X"d0",
X"0c",
X"ad",
X"f9",
X"07",
X"0d",
X"fa",
X"07",
X"d0",
X"04",
X"a9",
X"40",
X"85",
X"fc",
X"a9",
X"18",
X"8d",
X"87",
X"07",
X"a0",
X"23",
X"a9",
X"ff",
X"8d",
X"39",
X"01",
X"20",
X"5f",
X"8f",
X"a9",
X"a4",
X"4c",
X"06",
X"8f",
X"8d",
X"56",
X"07",
X"20",
X"31",
X"d9",
X"ee",
X"59",
X"07",
X"60",
X"ad",
X"23",
X"07",
X"f0",
X"fa",
X"a5",
X"ce",
X"25",
X"b5",
X"d0",
X"f4",
X"8d",
X"23",
X"07",
X"ee",
X"d6",
X"06",
X"4c",
X"98",
X"c9",
X"ad",
X"4e",
X"07",
X"d0",
X"37",
X"8d",
X"7d",
X"04",
X"ad",
X"47",
X"07",
X"d0",
X"2f",
X"a0",
X"04",
X"b9",
X"71",
X"04",
X"18",
X"79",
X"77",
X"04",
X"85",
X"02",
X"b9",
X"6b",
X"04",
X"f0",
X"1c",
X"69",
X"00",
X"85",
X"01",
X"a5",
X"86",
X"38",
X"f9",
X"71",
X"04",
X"a5",
X"6d",
X"f9",
X"6b",
X"04",
X"30",
X"0b",
X"a5",
X"02",
X"38",
X"e5",
X"86",
X"a5",
X"01",
X"e5",
X"6d",
X"10",
X"04",
X"88",
X"10",
X"d3",
X"60",
X"b9",
X"77",
X"04",
X"4a",
X"85",
X"00",
X"b9",
X"71",
X"04",
X"18",
X"65",
X"00",
X"85",
X"01",
X"b9",
X"6b",
X"04",
X"69",
X"00",
X"85",
X"00",
X"a5",
X"09",
X"4a",
X"90",
X"2c",
X"a5",
X"01",
X"38",
X"e5",
X"86",
X"a5",
X"00",
X"e5",
X"6d",
X"10",
X"0e",
X"a5",
X"86",
X"38",
X"e9",
X"01",
X"85",
X"86",
X"a5",
X"6d",
X"e9",
X"00",
X"4c",
X"39",
X"b8",
X"ad",
X"90",
X"04",
X"4a",
X"90",
X"0d",
X"a5",
X"86",
X"18",
X"69",
X"01",
X"85",
X"86",
X"a5",
X"6d",
X"69",
X"00",
X"85",
X"6d",
X"a9",
X"10",
X"85",
X"00",
X"a9",
X"01",
X"8d",
X"7d",
X"04",
X"85",
X"02",
X"4a",
X"aa",
X"4c",
X"d7",
X"bf",
X"05",
X"02",
X"08",
X"04",
X"01",
X"03",
X"03",
X"04",
X"04",
X"04",
X"a2",
X"05",
X"86",
X"08",
X"b5",
X"16",
X"c9",
X"30",
X"d0",
X"56",
X"a5",
X"0e",
X"c9",
X"04",
X"d0",
X"31",
X"a5",
X"1d",
X"c9",
X"03",
X"d0",
X"2b",
X"b5",
X"cf",
X"c9",
X"aa",
X"b0",
X"28",
X"a5",
X"ce",
X"c9",
X"a2",
X"b0",
X"22",
X"bd",
X"17",
X"04",
X"69",
X"ff",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"69",
X"01",
X"95",
X"cf",
X"ad",
X"0e",
X"01",
X"38",
X"e9",
X"ff",
X"8d",
X"0e",
X"01",
X"ad",
X"0d",
X"01",
X"e9",
X"01",
X"8d",
X"0d",
X"01",
X"4c",
X"ac",
X"b8",
X"ac",
X"0f",
X"01",
X"b9",
X"4b",
X"b8",
X"be",
X"50",
X"b8",
X"9d",
X"34",
X"01",
X"20",
X"27",
X"bc",
X"a9",
X"05",
X"85",
X"0e",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"4b",
X"e5",
X"60",
X"08",
X"10",
X"08",
X"00",
X"20",
X"af",
X"f1",
X"ad",
X"47",
X"07",
X"d0",
X"40",
X"ad",
X"0e",
X"07",
X"f0",
X"3b",
X"a8",
X"88",
X"98",
X"29",
X"02",
X"d0",
X"07",
X"e6",
X"ce",
X"e6",
X"ce",
X"4c",
X"d9",
X"b8",
X"c6",
X"ce",
X"c6",
X"ce",
X"b5",
X"58",
X"18",
X"79",
X"b6",
X"b8",
X"95",
X"cf",
X"c0",
X"01",
X"90",
X"0f",
X"a5",
X"0a",
X"29",
X"80",
X"f0",
X"09",
X"25",
X"0d",
X"d0",
X"05",
X"a9",
X"f4",
X"8d",
X"db",
X"06",
X"c0",
X"03",
X"d0",
X"0a",
X"ad",
X"db",
X"06",
X"85",
X"9f",
X"a9",
X"00",
X"8d",
X"0e",
X"07",
X"20",
X"52",
X"f1",
X"20",
X"7d",
X"e8",
X"20",
X"7a",
X"d6",
X"ad",
X"0e",
X"07",
X"f0",
X"0d",
X"ad",
X"86",
X"07",
X"d0",
X"08",
X"a9",
X"04",
X"8d",
X"86",
X"07",
X"ee",
X"0e",
X"07",
X"60",
X"a9",
X"2f",
X"95",
X"16",
X"a9",
X"01",
X"95",
X"0f",
X"b9",
X"76",
X"00",
X"95",
X"6e",
X"b9",
X"8f",
X"00",
X"95",
X"87",
X"b9",
X"d7",
X"00",
X"95",
X"cf",
X"ac",
X"98",
X"03",
X"d0",
X"03",
X"8d",
X"9d",
X"03",
X"8a",
X"99",
X"9a",
X"03",
X"ee",
X"98",
X"03",
X"a9",
X"04",
X"85",
X"fe",
X"60",
X"30",
X"60",
X"e0",
X"05",
X"d0",
X"68",
X"ac",
X"98",
X"03",
X"88",
X"ad",
X"99",
X"03",
X"d9",
X"49",
X"b9",
X"f0",
X"0f",
X"a5",
X"09",
X"4a",
X"4a",
X"90",
X"09",
X"a5",
X"d4",
X"e9",
X"01",
X"85",
X"d4",
X"ee",
X"99",
X"03",
X"ad",
X"99",
X"03",
X"c9",
X"08",
X"90",
X"46",
X"20",
X"52",
X"f1",
X"20",
X"af",
X"f1",
X"a0",
X"00",
X"20",
X"35",
X"e4",
X"c8",
X"cc",
X"98",
X"03",
X"d0",
X"f7",
X"ad",
X"d1",
X"03",
X"29",
X"0c",
X"f0",
X"10",
X"88",
X"be",
X"9a",
X"03",
X"20",
X"98",
X"c9",
X"88",
X"10",
X"f7",
X"8d",
X"98",
X"03",
X"8d",
X"99",
X"03",
X"ad",
X"99",
X"03",
X"c9",
X"20",
X"90",
X"17",
X"a2",
X"06",
X"a9",
X"01",
X"a0",
X"1b",
X"20",
X"f0",
X"e3",
X"a4",
X"02",
X"c0",
X"d0",
X"b0",
X"08",
X"b1",
X"06",
X"d0",
X"04",
X"a9",
X"26",
X"91",
X"06",
X"a6",
X"08",
X"60",
X"0f",
X"07",
X"ad",
X"4e",
X"07",
X"f0",
X"6f",
X"a2",
X"02",
X"86",
X"08",
X"b5",
X"0f",
X"d0",
X"51",
X"bd",
X"a8",
X"07",
X"ac",
X"cc",
X"06",
X"39",
X"ba",
X"b9",
X"c9",
X"06",
X"b0",
X"44",
X"a8",
X"b9",
X"6b",
X"04",
X"f0",
X"3e",
X"b9",
X"7d",
X"04",
X"f0",
X"08",
X"e9",
X"00",
X"99",
X"7d",
X"04",
X"4c",
X"1a",
X"ba",
X"ad",
X"47",
X"07",
X"d0",
X"2c",
X"a9",
X"0e",
X"99",
X"7d",
X"04",
X"b9",
X"6b",
X"04",
X"95",
X"6e",
X"b9",
X"71",
X"04",
X"95",
X"87",
X"b9",
X"77",
X"04",
X"38",
X"e9",
X"08",
X"95",
X"cf",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"4a",
X"95",
X"1e",
X"a9",
X"09",
X"9d",
X"9a",
X"04",
X"a9",
X"33",
X"95",
X"16",
X"4c",
X"2d",
X"ba",
X"b5",
X"16",
X"c9",
X"33",
X"d0",
X"0d",
X"20",
X"7a",
X"d6",
X"b5",
X"0f",
X"f0",
X"06",
X"20",
X"af",
X"f1",
X"20",
X"33",
X"ba",
X"ca",
X"10",
X"93",
X"60",
X"18",
X"e8",
X"ad",
X"47",
X"07",
X"d0",
X"3e",
X"b5",
X"1e",
X"d0",
X"2e",
X"ad",
X"d1",
X"03",
X"29",
X"0c",
X"c9",
X"0c",
X"f0",
X"40",
X"a0",
X"01",
X"20",
X"43",
X"e1",
X"30",
X"01",
X"c8",
X"94",
X"46",
X"88",
X"b9",
X"31",
X"ba",
X"95",
X"58",
X"a5",
X"00",
X"69",
X"28",
X"c9",
X"50",
X"90",
X"28",
X"a9",
X"01",
X"95",
X"1e",
X"a9",
X"0a",
X"9d",
X"8a",
X"07",
X"a9",
X"08",
X"85",
X"fe",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"03",
X"20",
X"63",
X"bf",
X"20",
X"02",
X"bf",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"43",
X"e2",
X"20",
X"53",
X"d8",
X"4c",
X"7d",
X"e8",
X"20",
X"98",
X"c9",
X"60",
X"04",
X"04",
X"04",
X"05",
X"05",
X"05",
X"06",
X"06",
X"06",
X"10",
X"f0",
X"ad",
X"a8",
X"07",
X"29",
X"07",
X"d0",
X"05",
X"ad",
X"a8",
X"07",
X"29",
X"08",
X"a8",
X"b9",
X"2a",
X"00",
X"d0",
X"19",
X"be",
X"89",
X"ba",
X"b5",
X"0f",
X"d0",
X"12",
X"a6",
X"08",
X"8a",
X"99",
X"ae",
X"06",
X"a9",
X"90",
X"99",
X"2a",
X"00",
X"a9",
X"07",
X"99",
X"a2",
X"04",
X"38",
X"60",
X"a6",
X"08",
X"18",
X"60",
X"ad",
X"47",
X"07",
X"d0",
X"63",
X"b5",
X"2a",
X"29",
X"7f",
X"bc",
X"ae",
X"06",
X"c9",
X"02",
X"f0",
X"20",
X"b0",
X"34",
X"8a",
X"18",
X"69",
X"0d",
X"aa",
X"a9",
X"10",
X"85",
X"00",
X"a9",
X"0f",
X"85",
X"01",
X"a9",
X"04",
X"85",
X"02",
X"a9",
X"00",
X"20",
X"d7",
X"bf",
X"20",
X"0f",
X"bf",
X"a6",
X"08",
X"4c",
X"28",
X"bb",
X"a9",
X"fe",
X"95",
X"ac",
X"b9",
X"1e",
X"00",
X"29",
X"f7",
X"99",
X"1e",
X"00",
X"b6",
X"46",
X"ca",
X"bd",
X"92",
X"ba",
X"a6",
X"08",
X"95",
X"64",
X"d6",
X"2a",
X"b9",
X"87",
X"00",
X"18",
X"69",
X"02",
X"95",
X"93",
X"b9",
X"6e",
X"00",
X"69",
X"00",
X"95",
X"7a",
X"b9",
X"cf",
X"00",
X"38",
X"e9",
X"0a",
X"95",
X"db",
X"a9",
X"01",
X"95",
X"c2",
X"d0",
X"03",
X"20",
X"c4",
X"d7",
X"20",
X"9b",
X"f1",
X"20",
X"48",
X"f1",
X"20",
X"36",
X"e2",
X"20",
X"dc",
X"e4",
X"60",
X"20",
X"84",
X"bb",
X"b5",
X"76",
X"99",
X"7a",
X"00",
X"b5",
X"8f",
X"09",
X"05",
X"99",
X"93",
X"00",
X"b5",
X"d7",
X"e9",
X"10",
X"99",
X"db",
X"00",
X"4c",
X"6c",
X"bb",
X"20",
X"84",
X"bb",
X"bd",
X"ea",
X"03",
X"99",
X"7a",
X"00",
X"a5",
X"06",
X"0a",
X"0a",
X"0a",
X"0a",
X"09",
X"05",
X"99",
X"93",
X"00",
X"a5",
X"02",
X"69",
X"20",
X"99",
X"db",
X"00",
X"a9",
X"fb",
X"99",
X"ac",
X"00",
X"a9",
X"01",
X"99",
X"c2",
X"00",
X"99",
X"2a",
X"00",
X"85",
X"fe",
X"86",
X"08",
X"20",
X"fe",
X"bb",
X"ee",
X"48",
X"07",
X"60",
X"a0",
X"08",
X"b9",
X"2a",
X"00",
X"f0",
X"07",
X"88",
X"c0",
X"05",
X"d0",
X"f6",
X"a0",
X"08",
X"8c",
X"b7",
X"06",
X"60",
X"a2",
X"08",
X"86",
X"08",
X"b5",
X"2a",
X"f0",
X"56",
X"0a",
X"90",
X"06",
X"20",
X"c3",
X"ba",
X"4c",
X"f4",
X"bb",
X"b4",
X"2a",
X"88",
X"f0",
X"1d",
X"f6",
X"2a",
X"b5",
X"93",
X"18",
X"6d",
X"75",
X"07",
X"95",
X"93",
X"b5",
X"7a",
X"69",
X"00",
X"95",
X"7a",
X"b5",
X"2a",
X"c9",
X"30",
X"d0",
X"26",
X"a9",
X"00",
X"95",
X"2a",
X"4c",
X"f4",
X"bb",
X"8a",
X"18",
X"69",
X"0d",
X"aa",
X"a9",
X"50",
X"85",
X"00",
X"a9",
X"06",
X"85",
X"02",
X"4a",
X"85",
X"01",
X"a9",
X"00",
X"20",
X"d7",
X"bf",
X"a6",
X"08",
X"b5",
X"ac",
X"c9",
X"05",
X"d0",
X"02",
X"f6",
X"2a",
X"20",
X"48",
X"f1",
X"20",
X"9b",
X"f1",
X"20",
X"36",
X"e2",
X"20",
X"86",
X"e6",
X"ca",
X"10",
X"a1",
X"60",
X"17",
X"1d",
X"0b",
X"11",
X"02",
X"13",
X"a9",
X"01",
X"8d",
X"39",
X"01",
X"ae",
X"53",
X"07",
X"bc",
X"f8",
X"bb",
X"20",
X"5f",
X"8f",
X"ee",
X"5e",
X"07",
X"ad",
X"5e",
X"07",
X"c9",
X"64",
X"d0",
X"0c",
X"a9",
X"00",
X"8d",
X"5e",
X"07",
X"ee",
X"5a",
X"07",
X"a9",
X"40",
X"85",
X"fe",
X"a9",
X"02",
X"8d",
X"38",
X"01",
X"ae",
X"53",
X"07",
X"bc",
X"fa",
X"bb",
X"20",
X"5f",
X"8f",
X"ac",
X"53",
X"07",
X"b9",
X"fc",
X"bb",
X"20",
X"06",
X"8f",
X"ac",
X"00",
X"03",
X"b9",
X"fb",
X"02",
X"d0",
X"05",
X"a9",
X"24",
X"99",
X"fb",
X"02",
X"a6",
X"08",
X"60",
X"a9",
X"2e",
X"85",
X"1b",
X"b5",
X"76",
X"85",
X"73",
X"b5",
X"8f",
X"85",
X"8c",
X"a9",
X"01",
X"85",
X"bb",
X"b5",
X"d7",
X"38",
X"e9",
X"08",
X"85",
X"d4",
X"a9",
X"01",
X"85",
X"23",
X"85",
X"14",
X"a9",
X"03",
X"8d",
X"9f",
X"04",
X"a5",
X"39",
X"c9",
X"02",
X"b0",
X"0a",
X"ad",
X"56",
X"07",
X"c9",
X"02",
X"90",
X"01",
X"4a",
X"85",
X"39",
X"a9",
X"20",
X"8d",
X"ca",
X"03",
X"a9",
X"02",
X"85",
X"fe",
X"60",
X"a2",
X"05",
X"86",
X"08",
X"a5",
X"23",
X"f0",
X"5d",
X"0a",
X"90",
X"23",
X"ad",
X"47",
X"07",
X"d0",
X"43",
X"a5",
X"39",
X"f0",
X"11",
X"c9",
X"03",
X"f0",
X"0d",
X"c9",
X"02",
X"d0",
X"37",
X"20",
X"f9",
X"ca",
X"20",
X"63",
X"e1",
X"4c",
X"d8",
X"bc",
X"20",
X"77",
X"ca",
X"20",
X"c1",
X"df",
X"4c",
X"d8",
X"bc",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"19",
X"c6",
X"d4",
X"a5",
X"23",
X"e6",
X"23",
X"c9",
X"11",
X"90",
X"0f",
X"a9",
X"10",
X"95",
X"58",
X"a9",
X"80",
X"85",
X"23",
X"0a",
X"8d",
X"ca",
X"03",
X"2a",
X"95",
X"46",
X"a5",
X"23",
X"c9",
X"06",
X"90",
X"12",
X"20",
X"52",
X"f1",
X"20",
X"af",
X"f1",
X"20",
X"43",
X"e2",
X"20",
X"d2",
X"e6",
X"20",
X"53",
X"d8",
X"20",
X"7a",
X"d6",
X"60",
X"04",
X"12",
X"48",
X"a9",
X"11",
X"ae",
X"ee",
X"03",
X"ac",
X"54",
X"07",
X"d0",
X"02",
X"a9",
X"12",
X"95",
X"26",
X"20",
X"6b",
X"8a",
X"ae",
X"ee",
X"03",
X"a5",
X"02",
X"9d",
X"e4",
X"03",
X"a8",
X"a5",
X"06",
X"9d",
X"e6",
X"03",
X"b1",
X"06",
X"20",
X"f6",
X"bd",
X"85",
X"00",
X"ac",
X"54",
X"07",
X"d0",
X"01",
X"98",
X"90",
X"25",
X"a0",
X"11",
X"94",
X"26",
X"a9",
X"c4",
X"a4",
X"00",
X"c0",
X"58",
X"f0",
X"04",
X"c0",
X"5d",
X"d0",
X"15",
X"ad",
X"bc",
X"06",
X"d0",
X"08",
X"a9",
X"0b",
X"8d",
X"9d",
X"07",
X"ee",
X"bc",
X"06",
X"ad",
X"9d",
X"07",
X"d0",
X"02",
X"a0",
X"c4",
X"98",
X"9d",
X"e8",
X"03",
X"20",
X"84",
X"bd",
X"a4",
X"02",
X"a9",
X"23",
X"91",
X"06",
X"a9",
X"10",
X"8d",
X"84",
X"07",
X"68",
X"85",
X"05",
X"a0",
X"00",
X"ad",
X"14",
X"07",
X"d0",
X"05",
X"ad",
X"54",
X"07",
X"f0",
X"01",
X"c8",
X"a5",
X"ce",
X"18",
X"79",
X"eb",
X"bc",
X"29",
X"f0",
X"95",
X"d7",
X"b4",
X"26",
X"c0",
X"11",
X"f0",
X"06",
X"20",
X"02",
X"be",
X"4c",
X"7b",
X"bd",
X"20",
X"9b",
X"bd",
X"ad",
X"ee",
X"03",
X"49",
X"01",
X"8d",
X"ee",
X"03",
X"60",
X"a5",
X"86",
X"18",
X"69",
X"08",
X"29",
X"f0",
X"95",
X"8f",
X"a5",
X"6d",
X"69",
X"00",
X"95",
X"76",
X"9d",
X"ea",
X"03",
X"a5",
X"b5",
X"95",
X"be",
X"60",
X"20",
X"1f",
X"be",
X"a9",
X"02",
X"85",
X"ff",
X"a9",
X"00",
X"95",
X"60",
X"9d",
X"3c",
X"04",
X"85",
X"9f",
X"a9",
X"fe",
X"95",
X"a8",
X"a5",
X"05",
X"20",
X"f6",
X"bd",
X"90",
X"31",
X"98",
X"c9",
X"09",
X"90",
X"02",
X"e9",
X"05",
X"20",
X"04",
X"8e",
X"d2",
X"bd",
X"38",
X"bb",
X"38",
X"bb",
X"d8",
X"bd",
X"d2",
X"bd",
X"df",
X"bd",
X"d5",
X"bd",
X"38",
X"bb",
X"d8",
X"bd",
X"a9",
X"00",
X"2c",
X"a9",
X"02",
X"2c",
X"a9",
X"03",
X"85",
X"39",
X"4c",
X"49",
X"bc",
X"a2",
X"05",
X"ac",
X"ee",
X"03",
X"20",
X"1e",
X"b9",
X"60",
X"c1",
X"c0",
X"5f",
X"60",
X"55",
X"56",
X"57",
X"58",
X"59",
X"5a",
X"5b",
X"5c",
X"5d",
X"5e",
X"a0",
X"0d",
X"d9",
X"e8",
X"bd",
X"f0",
X"04",
X"88",
X"10",
X"f8",
X"18",
X"60",
X"20",
X"1f",
X"be",
X"a9",
X"01",
X"9d",
X"ec",
X"03",
X"85",
X"fd",
X"20",
X"41",
X"be",
X"a9",
X"fe",
X"85",
X"9f",
X"a9",
X"05",
X"8d",
X"39",
X"01",
X"20",
X"27",
X"bc",
X"ae",
X"ee",
X"03",
X"60",
X"ae",
X"ee",
X"03",
X"a4",
X"02",
X"f0",
X"1a",
X"98",
X"38",
X"e9",
X"10",
X"85",
X"02",
X"a8",
X"b1",
X"06",
X"c9",
X"c2",
X"d0",
X"0d",
X"a9",
X"00",
X"91",
X"06",
X"20",
X"4d",
X"8a",
X"ae",
X"ee",
X"03",
X"20",
X"51",
X"bb",
X"60",
X"b5",
X"8f",
X"9d",
X"f1",
X"03",
X"a9",
X"f0",
X"95",
X"60",
X"95",
X"62",
X"a9",
X"fa",
X"95",
X"a8",
X"a9",
X"fc",
X"95",
X"aa",
X"a9",
X"00",
X"9d",
X"3c",
X"04",
X"9d",
X"3e",
X"04",
X"b5",
X"76",
X"95",
X"78",
X"b5",
X"8f",
X"95",
X"91",
X"b5",
X"d7",
X"18",
X"69",
X"08",
X"95",
X"d9",
X"a9",
X"fa",
X"95",
X"a8",
X"60",
X"b5",
X"26",
X"f0",
X"5d",
X"29",
X"0f",
X"48",
X"a8",
X"8a",
X"18",
X"69",
X"09",
X"aa",
X"88",
X"f0",
X"33",
X"20",
X"a4",
X"bf",
X"20",
X"0f",
X"bf",
X"8a",
X"18",
X"69",
X"02",
X"aa",
X"20",
X"a4",
X"bf",
X"20",
X"0f",
X"bf",
X"a6",
X"08",
X"20",
X"59",
X"f1",
X"20",
X"b6",
X"f1",
X"20",
X"53",
X"ec",
X"68",
X"b4",
X"be",
X"f0",
X"30",
X"48",
X"a9",
X"f0",
X"d5",
X"d9",
X"b0",
X"02",
X"95",
X"d9",
X"b5",
X"d7",
X"c9",
X"f0",
X"68",
X"90",
X"20",
X"b0",
X"1c",
X"20",
X"a4",
X"bf",
X"a6",
X"08",
X"20",
X"59",
X"f1",
X"20",
X"b6",
X"f1",
X"20",
X"d1",
X"eb",
X"b5",
X"d7",
X"29",
X"0f",
X"c9",
X"05",
X"68",
X"b0",
X"07",
X"a9",
X"01",
X"9d",
X"ec",
X"03",
X"a9",
X"00",
X"95",
X"26",
X"60",
X"a2",
X"01",
X"86",
X"08",
X"ad",
X"01",
X"03",
X"d0",
X"21",
X"bd",
X"ec",
X"03",
X"f0",
X"1c",
X"bd",
X"e6",
X"03",
X"85",
X"06",
X"a9",
X"05",
X"85",
X"07",
X"bd",
X"e4",
X"03",
X"85",
X"02",
X"a8",
X"bd",
X"e8",
X"03",
X"91",
X"06",
X"20",
X"61",
X"8a",
X"a9",
X"00",
X"9d",
X"ec",
X"03",
X"ca",
X"10",
X"d5",
X"60",
X"e8",
X"20",
X"0f",
X"bf",
X"a6",
X"08",
X"60",
X"ad",
X"0e",
X"07",
X"d0",
X"3e",
X"aa",
X"b5",
X"57",
X"0a",
X"0a",
X"0a",
X"0a",
X"85",
X"01",
X"b5",
X"57",
X"4a",
X"4a",
X"4a",
X"4a",
X"c9",
X"08",
X"90",
X"02",
X"09",
X"f0",
X"85",
X"00",
X"a0",
X"00",
X"c9",
X"00",
X"10",
X"01",
X"88",
X"84",
X"02",
X"bd",
X"00",
X"04",
X"18",
X"65",
X"01",
X"9d",
X"00",
X"04",
X"a9",
X"00",
X"2a",
X"48",
X"6a",
X"b5",
X"86",
X"65",
X"00",
X"95",
X"86",
X"b5",
X"6d",
X"65",
X"02",
X"95",
X"6d",
X"68",
X"18",
X"65",
X"00",
X"60",
X"a2",
X"00",
X"ad",
X"47",
X"07",
X"d0",
X"05",
X"ad",
X"0e",
X"07",
X"d0",
X"f3",
X"ad",
X"09",
X"07",
X"85",
X"00",
X"a9",
X"04",
X"4c",
X"ad",
X"bf",
X"a0",
X"3d",
X"b5",
X"1e",
X"c9",
X"05",
X"d0",
X"02",
X"a0",
X"20",
X"4c",
X"94",
X"bf",
X"a0",
X"00",
X"4c",
X"77",
X"bf",
X"a0",
X"01",
X"e8",
X"a9",
X"03",
X"85",
X"00",
X"a9",
X"06",
X"85",
X"01",
X"a9",
X"02",
X"85",
X"02",
X"98",
X"4c",
X"d1",
X"bf",
X"a0",
X"7f",
X"d0",
X"02",
X"a0",
X"0f",
X"a9",
X"02",
X"d0",
X"04",
X"a0",
X"1c",
X"a9",
X"03",
X"84",
X"00",
X"e8",
X"20",
X"ad",
X"bf",
X"a6",
X"08",
X"60",
X"06",
X"08",
X"a0",
X"00",
X"2c",
X"a0",
X"01",
X"a9",
X"50",
X"85",
X"00",
X"b9",
X"9f",
X"bf",
X"85",
X"02",
X"a9",
X"00",
X"4c",
X"d7",
X"bf",
X"a9",
X"00",
X"2c",
X"a9",
X"01",
X"48",
X"b4",
X"16",
X"e8",
X"a9",
X"05",
X"c0",
X"29",
X"d0",
X"02",
X"a9",
X"09",
X"85",
X"00",
X"a9",
X"0a",
X"85",
X"01",
X"a9",
X"03",
X"85",
X"02",
X"68",
X"a8",
X"20",
X"d7",
X"bf",
X"a6",
X"08",
X"60",
X"48",
X"bd",
X"16",
X"04",
X"18",
X"7d",
X"33",
X"04",
X"9d",
X"16",
X"04",
X"a0",
X"00",
X"b5",
X"9f",
X"10",
X"01",
X"88",
X"84",
X"07",
X"75",
X"ce",
X"95",
X"ce",
X"b5",
X"b5",
X"65",
X"07",
X"95",
X"b5",
X"bd",
X"33",
X"04",
X"18",
X"65",
X"00",
X"9d",
X"33",
X"04",
X"b5",
X"9f",
X"69",
X"00",
X"95",
X"9f",
X"c5",
X"02",
X"30",
X"10",
X"bd",
X"33",
X"04",
X"c9",
X"80",
X"90",
X"09",
X"a5",
X"02",
X"95",
X"9f",
X"a9",
X"00",
X"9d",
X"33",
X"04",
X"68",
X"f0",
X"2b",
X"a5",
X"02",
X"49",
X"ff",
X"a8",
X"c8",
X"84",
X"07",
X"bd",
X"33",
X"04",
X"38",
X"e5",
X"01",
X"9d",
X"33",
X"04",
X"b5",
X"9f",
X"e9",
X"00",
X"95",
X"9f",
X"c5",
X"07",
X"10",
X"10",
X"bd",
X"33",
X"04",
X"c9",
X"80",
X"b0",
X"09",
X"a5",
X"07",
X"95",
X"9f",
X"a9",
X"ff",
X"9d",
X"33",
X"04",
X"60",
X"b5",
X"0f",
X"48",
X"0a",
X"b0",
X"12",
X"68",
X"f0",
X"03",
X"4c",
X"82",
X"c8",
X"ad",
X"1f",
X"07",
X"29",
X"07",
X"c9",
X"07",
X"f0",
X"0e",
X"4c",
X"cc",
X"c0",
X"68",
X"29",
X"0f",
X"a8",
X"b9",
X"0f",
X"00",
X"d0",
X"02",
X"95",
X"0f",
X"60",
X"03",
X"03",
X"06",
X"06",
X"06",
X"06",
X"06",
X"06",
X"07",
X"07",
X"07",
X"05",
X"09",
X"04",
X"05",
X"06",
X"08",
X"09",
X"0a",
X"06",
X"0b",
X"10",
X"40",
X"b0",
X"b0",
X"80",
X"40",
X"40",
X"80",
X"40",
X"f0",
X"f0",
X"f0",
X"a5",
X"6d",
X"38",
X"e9",
X"04",
X"85",
X"6d",
X"ad",
X"25",
X"07",
X"38",
X"e9",
X"04",
X"8d",
X"25",
X"07",
X"ad",
X"1a",
X"07",
X"38",
X"e9",
X"04",
X"8d",
X"1a",
X"07",
X"ad",
X"1b",
X"07",
X"38",
X"e9",
X"04",
X"8d",
X"1b",
X"07",
X"ad",
X"2a",
X"07",
X"38",
X"e9",
X"04",
X"8d",
X"2a",
X"07",
X"a9",
X"00",
X"8d",
X"3b",
X"07",
X"8d",
X"2b",
X"07",
X"8d",
X"39",
X"07",
X"8d",
X"3a",
X"07",
X"b9",
X"f8",
X"9b",
X"8d",
X"2c",
X"07",
X"60",
X"ad",
X"45",
X"07",
X"f0",
X"5e",
X"ad",
X"26",
X"07",
X"d0",
X"59",
X"a0",
X"0b",
X"88",
X"30",
X"54",
X"ad",
X"5f",
X"07",
X"d9",
X"6b",
X"c0",
X"d0",
X"f5",
X"ad",
X"25",
X"07",
X"d9",
X"76",
X"c0",
X"d0",
X"ed",
X"a5",
X"ce",
X"d9",
X"81",
X"c0",
X"d0",
X"23",
X"a5",
X"1d",
X"c9",
X"00",
X"d0",
X"1d",
X"ad",
X"5f",
X"07",
X"c9",
X"06",
X"d0",
X"23",
X"ee",
X"d9",
X"06",
X"ee",
X"da",
X"06",
X"ad",
X"da",
X"06",
X"c9",
X"03",
X"d0",
X"1e",
X"ad",
X"d9",
X"06",
X"c9",
X"03",
X"f0",
X"0f",
X"d0",
X"07",
X"ad",
X"5f",
X"07",
X"c9",
X"06",
X"f0",
X"e6",
X"20",
X"8c",
X"c0",
X"20",
X"71",
X"d0",
X"a9",
X"00",
X"8d",
X"da",
X"06",
X"8d",
X"d9",
X"06",
X"a9",
X"00",
X"8d",
X"45",
X"07",
X"ad",
X"cd",
X"06",
X"f0",
X"10",
X"95",
X"16",
X"a9",
X"01",
X"95",
X"0f",
X"a9",
X"00",
X"95",
X"1e",
X"8d",
X"cd",
X"06",
X"4c",
X"26",
X"c2",
X"ac",
X"39",
X"07",
X"b1",
X"e9",
X"c9",
X"ff",
X"d0",
X"03",
X"4c",
X"16",
X"c2",
X"29",
X"0f",
X"c9",
X"0e",
X"f0",
X"0e",
X"e0",
X"05",
X"90",
X"0a",
X"c8",
X"b1",
X"e9",
X"29",
X"3f",
X"c9",
X"2e",
X"f0",
X"01",
X"60",
X"ad",
X"1d",
X"07",
X"18",
X"69",
X"30",
X"29",
X"f0",
X"85",
X"07",
X"ad",
X"1b",
X"07",
X"69",
X"00",
X"85",
X"06",
X"ac",
X"39",
X"07",
X"c8",
X"b1",
X"e9",
X"0a",
X"90",
X"0b",
X"ad",
X"3b",
X"07",
X"d0",
X"06",
X"ee",
X"3b",
X"07",
X"ee",
X"3a",
X"07",
X"88",
X"b1",
X"e9",
X"29",
X"0f",
X"c9",
X"0f",
X"d0",
X"19",
X"ad",
X"3b",
X"07",
X"d0",
X"14",
X"c8",
X"b1",
X"e9",
X"29",
X"3f",
X"8d",
X"3a",
X"07",
X"ee",
X"39",
X"07",
X"ee",
X"39",
X"07",
X"ee",
X"3b",
X"07",
X"4c",
X"cc",
X"c0",
X"ad",
X"3a",
X"07",
X"95",
X"6e",
X"b1",
X"e9",
X"29",
X"f0",
X"95",
X"87",
X"cd",
X"1d",
X"07",
X"b5",
X"6e",
X"ed",
X"1b",
X"07",
X"b0",
X"0b",
X"b1",
X"e9",
X"29",
X"0f",
X"c9",
X"0e",
X"f0",
X"69",
X"4c",
X"50",
X"c2",
X"a5",
X"07",
X"d5",
X"87",
X"a5",
X"06",
X"f5",
X"6e",
X"90",
X"41",
X"a9",
X"01",
X"95",
X"b6",
X"b1",
X"e9",
X"0a",
X"0a",
X"0a",
X"0a",
X"95",
X"cf",
X"c9",
X"e0",
X"f0",
X"4c",
X"c8",
X"b1",
X"e9",
X"29",
X"40",
X"f0",
X"05",
X"ad",
X"cc",
X"06",
X"f0",
X"6d",
X"b1",
X"e9",
X"29",
X"3f",
X"c9",
X"37",
X"90",
X"04",
X"c9",
X"3f",
X"90",
X"31",
X"c9",
X"06",
X"d0",
X"07",
X"ac",
X"6a",
X"07",
X"f0",
X"02",
X"a9",
X"02",
X"95",
X"16",
X"a9",
X"01",
X"95",
X"0f",
X"20",
X"26",
X"c2",
X"b5",
X"0f",
X"d0",
X"49",
X"60",
X"ad",
X"cb",
X"06",
X"d0",
X"09",
X"ad",
X"98",
X"03",
X"c9",
X"01",
X"d0",
X"0b",
X"a9",
X"2f",
X"95",
X"16",
X"a9",
X"00",
X"95",
X"1e",
X"20",
X"6c",
X"c2",
X"60",
X"4c",
X"1b",
X"c7",
X"c8",
X"c8",
X"b1",
X"e9",
X"4a",
X"4a",
X"4a",
X"4a",
X"4a",
X"cd",
X"5f",
X"07",
X"d0",
X"0e",
X"88",
X"b1",
X"e9",
X"8d",
X"50",
X"07",
X"c8",
X"b1",
X"e9",
X"29",
X"1f",
X"8d",
X"51",
X"07",
X"4c",
X"5b",
X"c2",
X"ac",
X"39",
X"07",
X"b1",
X"e9",
X"29",
X"0f",
X"c9",
X"0e",
X"d0",
X"03",
X"ee",
X"39",
X"07",
X"ee",
X"39",
X"07",
X"ee",
X"39",
X"07",
X"a9",
X"00",
X"8d",
X"3b",
X"07",
X"a6",
X"08",
X"60",
X"b5",
X"16",
X"c9",
X"15",
X"b0",
X"0d",
X"a8",
X"b5",
X"cf",
X"69",
X"08",
X"95",
X"cf",
X"a9",
X"01",
X"9d",
X"d8",
X"03",
X"98",
X"20",
X"04",
X"8e",
X"0e",
X"c3",
X"0e",
X"c3",
X"0e",
X"c3",
X"1e",
X"c3",
X"f0",
X"c2",
X"28",
X"c3",
X"f1",
X"c2",
X"42",
X"c3",
X"6b",
X"c3",
X"f0",
X"c2",
X"75",
X"c3",
X"75",
X"c3",
X"f7",
X"c2",
X"87",
X"c7",
X"d1",
X"c7",
X"4a",
X"c3",
X"3d",
X"c3",
X"85",
X"c3",
X"a0",
X"c7",
X"f0",
X"c2",
X"a0",
X"c7",
X"a0",
X"c7",
X"a0",
X"c7",
X"a0",
X"c7",
X"b8",
X"c7",
X"f0",
X"c2",
X"f0",
X"c2",
X"5c",
X"c4",
X"5c",
X"c4",
X"5c",
X"c4",
X"5c",
X"c4",
X"59",
X"c4",
X"f0",
X"c2",
X"f0",
X"c2",
X"f0",
X"c2",
X"f0",
X"c2",
X"df",
X"c7",
X"12",
X"c8",
X"3f",
X"c8",
X"45",
X"c8",
X"0b",
X"c8",
X"03",
X"c8",
X"0b",
X"c8",
X"4b",
X"c8",
X"57",
X"c8",
X"49",
X"c5",
X"60",
X"bc",
X"1e",
X"b9",
X"f0",
X"c2",
X"f0",
X"c2",
X"f0",
X"c2",
X"f0",
X"c2",
X"f0",
X"c2",
X"07",
X"c3",
X"81",
X"c8",
X"60",
X"20",
X"0e",
X"c3",
X"4c",
X"46",
X"c3",
X"a9",
X"02",
X"95",
X"b6",
X"95",
X"cf",
X"4a",
X"9d",
X"96",
X"07",
X"4a",
X"95",
X"1e",
X"4c",
X"46",
X"c3",
X"a9",
X"b8",
X"95",
X"cf",
X"60",
X"f8",
X"f4",
X"a0",
X"01",
X"ad",
X"6a",
X"07",
X"d0",
X"01",
X"88",
X"b9",
X"0c",
X"c3",
X"95",
X"58",
X"4c",
X"5a",
X"c3",
X"20",
X"0e",
X"c3",
X"a9",
X"01",
X"95",
X"1e",
X"60",
X"80",
X"50",
X"a9",
X"00",
X"9d",
X"a2",
X"03",
X"95",
X"58",
X"ac",
X"cc",
X"06",
X"b9",
X"26",
X"c3",
X"9d",
X"96",
X"07",
X"a9",
X"0b",
X"4c",
X"5c",
X"c3",
X"a9",
X"00",
X"4c",
X"19",
X"c3",
X"a9",
X"00",
X"95",
X"58",
X"a9",
X"09",
X"d0",
X"12",
X"a0",
X"30",
X"b5",
X"cf",
X"9d",
X"01",
X"04",
X"10",
X"02",
X"a0",
X"e0",
X"98",
X"75",
X"cf",
X"95",
X"58",
X"a9",
X"03",
X"9d",
X"9a",
X"04",
X"a9",
X"02",
X"95",
X"46",
X"a9",
X"00",
X"95",
X"a0",
X"9d",
X"34",
X"04",
X"60",
X"a9",
X"02",
X"95",
X"46",
X"a9",
X"09",
X"9d",
X"9a",
X"04",
X"60",
X"20",
X"46",
X"c3",
X"bd",
X"a7",
X"07",
X"29",
X"10",
X"95",
X"58",
X"b5",
X"cf",
X"9d",
X"34",
X"04",
X"60",
X"ad",
X"cb",
X"06",
X"d0",
X"0b",
X"a9",
X"00",
X"8d",
X"d1",
X"06",
X"20",
X"3d",
X"c3",
X"4c",
X"d9",
X"c7",
X"4c",
X"98",
X"c9",
X"26",
X"2c",
X"32",
X"38",
X"20",
X"22",
X"24",
X"26",
X"13",
X"14",
X"15",
X"16",
X"ad",
X"8f",
X"07",
X"d0",
X"3c",
X"e0",
X"05",
X"b0",
X"38",
X"a9",
X"80",
X"8d",
X"8f",
X"07",
X"a0",
X"04",
X"b9",
X"16",
X"00",
X"c9",
X"11",
X"f0",
X"2b",
X"88",
X"10",
X"f6",
X"ee",
X"d1",
X"06",
X"ad",
X"d1",
X"06",
X"c9",
X"07",
X"90",
X"1d",
X"a2",
X"04",
X"b5",
X"0f",
X"f0",
X"05",
X"ca",
X"10",
X"f9",
X"30",
X"10",
X"a9",
X"00",
X"95",
X"1e",
X"a9",
X"11",
X"95",
X"16",
X"20",
X"8a",
X"c3",
X"a9",
X"20",
X"20",
X"d8",
X"c5",
X"a6",
X"08",
X"60",
X"a5",
X"ce",
X"c9",
X"2c",
X"90",
X"f9",
X"b9",
X"1e",
X"00",
X"d0",
X"f4",
X"b9",
X"6e",
X"00",
X"95",
X"6e",
X"b9",
X"87",
X"00",
X"95",
X"87",
X"a9",
X"01",
X"95",
X"b6",
X"b9",
X"cf",
X"00",
X"38",
X"e9",
X"08",
X"95",
X"cf",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"a8",
X"a2",
X"02",
X"b9",
X"98",
X"c3",
X"95",
X"01",
X"c8",
X"c8",
X"c8",
X"c8",
X"ca",
X"10",
X"f4",
X"a6",
X"08",
X"20",
X"6c",
X"cf",
X"a4",
X"57",
X"c0",
X"08",
X"b0",
X"0e",
X"a8",
X"bd",
X"a8",
X"07",
X"29",
X"03",
X"f0",
X"05",
X"98",
X"49",
X"ff",
X"a8",
X"c8",
X"98",
X"20",
X"46",
X"c3",
X"a0",
X"02",
X"95",
X"58",
X"c9",
X"00",
X"30",
X"01",
X"88",
X"94",
X"46",
X"a9",
X"fd",
X"95",
X"a0",
X"a9",
X"01",
X"95",
X"0f",
X"a9",
X"05",
X"95",
X"1e",
X"60",
X"28",
X"38",
X"28",
X"38",
X"28",
X"00",
X"00",
X"10",
X"10",
X"00",
X"20",
X"75",
X"c5",
X"a9",
X"00",
X"95",
X"58",
X"b5",
X"16",
X"38",
X"e9",
X"1b",
X"a8",
X"b9",
X"4f",
X"c4",
X"9d",
X"88",
X"03",
X"b9",
X"54",
X"c4",
X"95",
X"34",
X"b5",
X"cf",
X"18",
X"69",
X"04",
X"95",
X"cf",
X"b5",
X"87",
X"18",
X"69",
X"04",
X"95",
X"87",
X"b5",
X"6e",
X"69",
X"00",
X"95",
X"6e",
X"4c",
X"d9",
X"c7",
X"80",
X"30",
X"40",
X"80",
X"30",
X"50",
X"50",
X"70",
X"20",
X"40",
X"80",
X"a0",
X"70",
X"40",
X"90",
X"68",
X"0e",
X"05",
X"06",
X"0e",
X"1c",
X"20",
X"10",
X"0c",
X"1e",
X"22",
X"18",
X"14",
X"10",
X"60",
X"20",
X"48",
X"ad",
X"8f",
X"07",
X"d0",
X"a1",
X"20",
X"46",
X"c3",
X"bd",
X"a8",
X"07",
X"29",
X"03",
X"a8",
X"b9",
X"a4",
X"c4",
X"8d",
X"8f",
X"07",
X"a0",
X"03",
X"ad",
X"cc",
X"06",
X"f0",
X"01",
X"c8",
X"84",
X"00",
X"e4",
X"00",
X"b0",
X"84",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"85",
X"00",
X"85",
X"01",
X"a9",
X"fb",
X"95",
X"a0",
X"a9",
X"00",
X"a4",
X"57",
X"f0",
X"07",
X"a9",
X"04",
X"c0",
X"19",
X"90",
X"01",
X"0a",
X"48",
X"18",
X"65",
X"00",
X"85",
X"00",
X"bd",
X"a8",
X"07",
X"29",
X"03",
X"f0",
X"07",
X"bd",
X"a9",
X"07",
X"29",
X"0f",
X"85",
X"00",
X"68",
X"18",
X"65",
X"01",
X"a8",
X"b9",
X"98",
X"c4",
X"95",
X"58",
X"a9",
X"01",
X"95",
X"46",
X"a5",
X"57",
X"d0",
X"12",
X"a4",
X"00",
X"98",
X"29",
X"02",
X"f0",
X"0b",
X"b5",
X"58",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"95",
X"58",
X"f6",
X"46",
X"98",
X"29",
X"02",
X"f0",
X"0f",
X"a5",
X"86",
X"18",
X"79",
X"88",
X"c4",
X"95",
X"87",
X"a5",
X"6d",
X"69",
X"00",
X"4c",
X"3c",
X"c5",
X"a5",
X"86",
X"38",
X"f9",
X"88",
X"c4",
X"95",
X"87",
X"a5",
X"6d",
X"e9",
X"00",
X"95",
X"6e",
X"a9",
X"01",
X"95",
X"0f",
X"95",
X"b6",
X"a9",
X"f8",
X"95",
X"cf",
X"60",
X"20",
X"75",
X"c5",
X"8e",
X"68",
X"03",
X"a9",
X"00",
X"8d",
X"63",
X"03",
X"8d",
X"69",
X"03",
X"b5",
X"87",
X"8d",
X"66",
X"03",
X"a9",
X"df",
X"8d",
X"90",
X"07",
X"95",
X"46",
X"a9",
X"20",
X"8d",
X"64",
X"03",
X"9d",
X"8a",
X"07",
X"a9",
X"05",
X"8d",
X"83",
X"04",
X"4a",
X"8d",
X"65",
X"03",
X"60",
X"a0",
X"ff",
X"c8",
X"b9",
X"0f",
X"00",
X"d0",
X"fa",
X"8c",
X"cf",
X"06",
X"8a",
X"09",
X"80",
X"99",
X"0f",
X"00",
X"b5",
X"6e",
X"99",
X"6e",
X"00",
X"b5",
X"87",
X"99",
X"87",
X"00",
X"a9",
X"01",
X"95",
X"0f",
X"99",
X"b6",
X"00",
X"b5",
X"cf",
X"99",
X"cf",
X"00",
X"60",
X"90",
X"80",
X"70",
X"90",
X"ff",
X"01",
X"ad",
X"8f",
X"07",
X"d0",
X"f4",
X"9d",
X"34",
X"04",
X"a5",
X"fd",
X"09",
X"02",
X"85",
X"fd",
X"ac",
X"68",
X"03",
X"b9",
X"16",
X"00",
X"c9",
X"2d",
X"f0",
X"31",
X"20",
X"d9",
X"d1",
X"18",
X"69",
X"20",
X"ac",
X"cc",
X"06",
X"f0",
X"03",
X"38",
X"e9",
X"10",
X"8d",
X"8f",
X"07",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"9d",
X"17",
X"04",
X"a8",
X"b9",
X"9d",
X"c5",
X"95",
X"cf",
X"ad",
X"1d",
X"07",
X"18",
X"69",
X"20",
X"95",
X"87",
X"ad",
X"1b",
X"07",
X"69",
X"00",
X"95",
X"6e",
X"4c",
X"1f",
X"c6",
X"b9",
X"87",
X"00",
X"38",
X"e9",
X"0e",
X"95",
X"87",
X"b9",
X"6e",
X"00",
X"95",
X"6e",
X"b9",
X"cf",
X"00",
X"18",
X"69",
X"08",
X"95",
X"cf",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"9d",
X"17",
X"04",
X"a8",
X"b9",
X"9d",
X"c5",
X"a0",
X"00",
X"d5",
X"cf",
X"90",
X"01",
X"c8",
X"b9",
X"a1",
X"c5",
X"9d",
X"34",
X"04",
X"a9",
X"00",
X"8d",
X"cb",
X"06",
X"a9",
X"08",
X"9d",
X"9a",
X"04",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"4a",
X"9d",
X"01",
X"04",
X"95",
X"1e",
X"60",
X"00",
X"30",
X"60",
X"60",
X"00",
X"20",
X"60",
X"40",
X"70",
X"40",
X"60",
X"30",
X"ad",
X"8f",
X"07",
X"d0",
X"47",
X"a9",
X"20",
X"8d",
X"8f",
X"07",
X"ce",
X"d7",
X"06",
X"a0",
X"06",
X"88",
X"b9",
X"16",
X"00",
X"c9",
X"31",
X"d0",
X"f8",
X"b9",
X"87",
X"00",
X"38",
X"e9",
X"30",
X"48",
X"b9",
X"6e",
X"00",
X"e9",
X"00",
X"85",
X"00",
X"ad",
X"d7",
X"06",
X"18",
X"79",
X"1e",
X"00",
X"a8",
X"68",
X"18",
X"79",
X"31",
X"c6",
X"95",
X"87",
X"a5",
X"00",
X"69",
X"00",
X"95",
X"6e",
X"b9",
X"37",
X"c6",
X"95",
X"cf",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"4a",
X"95",
X"58",
X"a9",
X"08",
X"95",
X"a0",
X"60",
X"01",
X"02",
X"04",
X"08",
X"10",
X"20",
X"40",
X"80",
X"40",
X"30",
X"90",
X"50",
X"20",
X"60",
X"a0",
X"70",
X"0a",
X"0b",
X"ad",
X"8f",
X"07",
X"d0",
X"6f",
X"ad",
X"4e",
X"07",
X"d0",
X"57",
X"e0",
X"03",
X"b0",
X"66",
X"a0",
X"00",
X"bd",
X"a7",
X"07",
X"c9",
X"aa",
X"90",
X"01",
X"c8",
X"ad",
X"5f",
X"07",
X"c9",
X"01",
X"f0",
X"01",
X"c8",
X"98",
X"29",
X"01",
X"a8",
X"b9",
X"9a",
X"c6",
X"95",
X"16",
X"ad",
X"dd",
X"06",
X"c9",
X"ff",
X"d0",
X"05",
X"a9",
X"00",
X"8d",
X"dd",
X"06",
X"bd",
X"a7",
X"07",
X"29",
X"07",
X"a8",
X"b9",
X"8a",
X"c6",
X"2c",
X"dd",
X"06",
X"f0",
X"07",
X"c8",
X"98",
X"29",
X"07",
X"4c",
X"d6",
X"c6",
X"0d",
X"dd",
X"06",
X"8d",
X"dd",
X"06",
X"b9",
X"92",
X"c6",
X"20",
X"d8",
X"c5",
X"9d",
X"17",
X"04",
X"a9",
X"20",
X"8d",
X"8f",
X"07",
X"4c",
X"6c",
X"c2",
X"a0",
X"ff",
X"c8",
X"c0",
X"05",
X"b0",
X"0d",
X"b9",
X"0f",
X"00",
X"f0",
X"f6",
X"b9",
X"16",
X"00",
X"c9",
X"08",
X"d0",
X"ef",
X"60",
X"a5",
X"fe",
X"09",
X"08",
X"85",
X"fe",
X"a9",
X"08",
X"d0",
X"a8",
X"a0",
X"00",
X"38",
X"e9",
X"37",
X"48",
X"c9",
X"04",
X"b0",
X"0b",
X"48",
X"a0",
X"06",
X"ad",
X"6a",
X"07",
X"f0",
X"02",
X"a0",
X"02",
X"68",
X"84",
X"01",
X"a0",
X"b0",
X"29",
X"02",
X"f0",
X"02",
X"a0",
X"70",
X"84",
X"00",
X"ad",
X"1b",
X"07",
X"85",
X"02",
X"ad",
X"1d",
X"07",
X"85",
X"03",
X"a0",
X"02",
X"68",
X"4a",
X"90",
X"01",
X"c8",
X"8c",
X"d3",
X"06",
X"a2",
X"ff",
X"e8",
X"e0",
X"05",
X"b0",
X"2d",
X"b5",
X"0f",
X"d0",
X"f7",
X"a5",
X"01",
X"95",
X"16",
X"a5",
X"02",
X"95",
X"6e",
X"a5",
X"03",
X"95",
X"87",
X"18",
X"69",
X"18",
X"85",
X"03",
X"a5",
X"02",
X"69",
X"00",
X"85",
X"02",
X"a5",
X"00",
X"95",
X"cf",
X"a9",
X"01",
X"95",
X"b6",
X"95",
X"0f",
X"20",
X"6c",
X"c2",
X"ce",
X"d3",
X"06",
X"d0",
X"cc",
X"4c",
X"5e",
X"c2",
X"a9",
X"01",
X"95",
X"58",
X"4a",
X"95",
X"1e",
X"95",
X"a0",
X"b5",
X"cf",
X"9d",
X"34",
X"04",
X"38",
X"e9",
X"18",
X"9d",
X"17",
X"04",
X"a9",
X"09",
X"4c",
X"db",
X"c7",
X"b5",
X"16",
X"8d",
X"cb",
X"06",
X"38",
X"e9",
X"12",
X"20",
X"04",
X"8e",
X"a4",
X"c3",
X"b7",
X"c7",
X"a8",
X"c4",
X"a3",
X"c5",
X"3d",
X"c6",
X"9c",
X"c6",
X"60",
X"a0",
X"05",
X"b9",
X"16",
X"00",
X"c9",
X"11",
X"d0",
X"05",
X"a9",
X"01",
X"99",
X"1e",
X"00",
X"88",
X"10",
X"f1",
X"a9",
X"00",
X"8d",
X"cb",
X"06",
X"95",
X"0f",
X"60",
X"a9",
X"02",
X"95",
X"46",
X"a9",
X"f8",
X"95",
X"58",
X"a9",
X"03",
X"9d",
X"9a",
X"04",
X"60",
X"d6",
X"cf",
X"d6",
X"cf",
X"ac",
X"cc",
X"06",
X"d0",
X"05",
X"a0",
X"02",
X"20",
X"71",
X"c8",
X"a0",
X"ff",
X"ad",
X"a0",
X"03",
X"95",
X"1e",
X"10",
X"02",
X"8a",
X"a8",
X"8c",
X"a0",
X"03",
X"a9",
X"00",
X"95",
X"46",
X"a8",
X"20",
X"71",
X"c8",
X"a9",
X"ff",
X"9d",
X"a2",
X"03",
X"4c",
X"28",
X"c8",
X"a9",
X"00",
X"95",
X"58",
X"4c",
X"28",
X"c8",
X"a0",
X"40",
X"b5",
X"cf",
X"10",
X"07",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"a0",
X"c0",
X"9d",
X"01",
X"04",
X"98",
X"18",
X"75",
X"cf",
X"95",
X"58",
X"20",
X"63",
X"c3",
X"a9",
X"05",
X"ac",
X"4e",
X"07",
X"c0",
X"03",
X"f0",
X"07",
X"ac",
X"cc",
X"06",
X"d0",
X"02",
X"a9",
X"06",
X"9d",
X"9a",
X"04",
X"60",
X"20",
X"4b",
X"c8",
X"4c",
X"48",
X"c8",
X"20",
X"57",
X"c8",
X"4c",
X"2b",
X"c8",
X"a9",
X"10",
X"9d",
X"34",
X"04",
X"a9",
X"ff",
X"95",
X"a0",
X"4c",
X"60",
X"c8",
X"a9",
X"f0",
X"9d",
X"34",
X"04",
X"a9",
X"00",
X"95",
X"a0",
X"a0",
X"01",
X"20",
X"71",
X"c8",
X"a9",
X"04",
X"9d",
X"9a",
X"04",
X"60",
X"08",
X"0c",
X"f8",
X"00",
X"00",
X"ff",
X"b5",
X"87",
X"18",
X"79",
X"6b",
X"c8",
X"95",
X"87",
X"b5",
X"6e",
X"79",
X"6e",
X"c8",
X"95",
X"6e",
X"60",
X"60",
X"a6",
X"08",
X"a9",
X"00",
X"b4",
X"16",
X"c0",
X"15",
X"90",
X"03",
X"98",
X"e9",
X"14",
X"20",
X"04",
X"8e",
X"e0",
X"c8",
X"35",
X"c9",
X"95",
X"d2",
X"d6",
X"c8",
X"d6",
X"c8",
X"d6",
X"c8",
X"d6",
X"c8",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"47",
X"c9",
X"d6",
X"c8",
X"65",
X"c9",
X"65",
X"c9",
X"65",
X"c9",
X"65",
X"c9",
X"65",
X"c9",
X"65",
X"c9",
X"65",
X"c9",
X"4d",
X"c9",
X"4d",
X"c9",
X"65",
X"d0",
X"85",
X"bc",
X"4b",
X"b9",
X"d6",
X"c8",
X"d9",
X"d2",
X"ba",
X"b8",
X"d6",
X"c8",
X"a4",
X"b7",
X"d7",
X"c8",
X"60",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"4c",
X"7d",
X"e8",
X"a9",
X"00",
X"9d",
X"c5",
X"03",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"7d",
X"e8",
X"20",
X"43",
X"e2",
X"20",
X"c1",
X"df",
X"20",
X"33",
X"da",
X"20",
X"53",
X"d8",
X"ac",
X"47",
X"07",
X"d0",
X"03",
X"20",
X"05",
X"c9",
X"4c",
X"7a",
X"d6",
X"b5",
X"16",
X"20",
X"04",
X"8e",
X"77",
X"ca",
X"77",
X"ca",
X"77",
X"ca",
X"77",
X"ca",
X"77",
X"ca",
X"d8",
X"c9",
X"77",
X"ca",
X"89",
X"cb",
X"36",
X"cc",
X"34",
X"c9",
X"4a",
X"cc",
X"4a",
X"cc",
X"b0",
X"c9",
X"b0",
X"d3",
X"f9",
X"ca",
X"ff",
X"ca",
X"25",
X"cb",
X"28",
X"cf",
X"77",
X"ca",
X"34",
X"c9",
X"df",
X"ce",
X"60",
X"20",
X"eb",
X"d1",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"43",
X"e2",
X"20",
X"53",
X"d8",
X"4c",
X"7a",
X"d6",
X"20",
X"3c",
X"cd",
X"4c",
X"7a",
X"d6",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"4c",
X"e2",
X"20",
X"7b",
X"db",
X"20",
X"52",
X"f1",
X"20",
X"66",
X"ed",
X"20",
X"55",
X"d6",
X"4c",
X"7a",
X"d6",
X"20",
X"af",
X"f1",
X"20",
X"52",
X"f1",
X"20",
X"73",
X"e2",
X"20",
X"45",
X"db",
X"ad",
X"47",
X"07",
X"d0",
X"03",
X"20",
X"82",
X"c9",
X"20",
X"52",
X"f1",
X"20",
X"c8",
X"e5",
X"4c",
X"7a",
X"d6",
X"b5",
X"16",
X"38",
X"e9",
X"24",
X"20",
X"04",
X"8e",
X"32",
X"d4",
X"d3",
X"d5",
X"4f",
X"d6",
X"4f",
X"d6",
X"07",
X"d6",
X"31",
X"d6",
X"3d",
X"d6",
X"a9",
X"00",
X"95",
X"0f",
X"95",
X"16",
X"95",
X"1e",
X"9d",
X"10",
X"01",
X"9d",
X"96",
X"07",
X"9d",
X"25",
X"01",
X"9d",
X"c5",
X"03",
X"9d",
X"8a",
X"07",
X"60",
X"bd",
X"96",
X"07",
X"d0",
X"16",
X"20",
X"f7",
X"c2",
X"bd",
X"a8",
X"07",
X"09",
X"80",
X"9d",
X"34",
X"04",
X"29",
X"0f",
X"09",
X"06",
X"9d",
X"96",
X"07",
X"a9",
X"f9",
X"95",
X"a0",
X"4c",
X"92",
X"bf",
X"30",
X"1c",
X"00",
X"e8",
X"00",
X"18",
X"08",
X"f8",
X"0c",
X"f4",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"03",
X"4c",
X"e5",
X"ca",
X"b5",
X"3c",
X"f0",
X"2d",
X"d6",
X"3c",
X"ad",
X"d1",
X"03",
X"29",
X"0c",
X"d0",
X"6a",
X"bd",
X"a2",
X"03",
X"d0",
X"17",
X"ac",
X"cc",
X"06",
X"b9",
X"ce",
X"c9",
X"9d",
X"a2",
X"03",
X"20",
X"94",
X"ba",
X"90",
X"09",
X"b5",
X"1e",
X"09",
X"08",
X"95",
X"1e",
X"4c",
X"58",
X"ca",
X"de",
X"a2",
X"03",
X"4c",
X"58",
X"ca",
X"20",
X"37",
X"b5",
X"1e",
X"29",
X"07",
X"c9",
X"01",
X"f0",
X"3e",
X"a9",
X"00",
X"85",
X"00",
X"a0",
X"fa",
X"b5",
X"cf",
X"30",
X"13",
X"a0",
X"fd",
X"c9",
X"70",
X"e6",
X"00",
X"90",
X"0b",
X"c6",
X"00",
X"bd",
X"a8",
X"07",
X"29",
X"01",
X"d0",
X"02",
X"a0",
X"fa",
X"94",
X"a0",
X"b5",
X"1e",
X"09",
X"01",
X"95",
X"1e",
X"a5",
X"00",
X"3d",
X"a9",
X"07",
X"a8",
X"ad",
X"cc",
X"06",
X"d0",
X"01",
X"a8",
X"b9",
X"10",
X"ca",
X"9d",
X"8a",
X"07",
X"bd",
X"a8",
X"07",
X"09",
X"c0",
X"95",
X"3c",
X"a0",
X"fc",
X"a5",
X"09",
X"29",
X"40",
X"d0",
X"02",
X"a0",
X"04",
X"94",
X"58",
X"a0",
X"01",
X"20",
X"43",
X"e1",
X"30",
X"0a",
X"c8",
X"bd",
X"96",
X"07",
X"d0",
X"04",
X"a9",
X"f8",
X"95",
X"58",
X"94",
X"46",
X"a0",
X"00",
X"b5",
X"1e",
X"29",
X"40",
X"d0",
X"19",
X"b5",
X"1e",
X"0a",
X"b0",
X"30",
X"b5",
X"1e",
X"29",
X"20",
X"d0",
X"5b",
X"b5",
X"1e",
X"29",
X"07",
X"f0",
X"24",
X"c9",
X"05",
X"f0",
X"04",
X"c9",
X"03",
X"b0",
X"30",
X"20",
X"63",
X"bf",
X"a0",
X"00",
X"b5",
X"1e",
X"c9",
X"02",
X"f0",
X"0c",
X"29",
X"40",
X"f0",
X"0d",
X"b5",
X"16",
X"c9",
X"2e",
X"f0",
X"07",
X"d0",
X"03",
X"4c",
X"02",
X"bf",
X"a0",
X"01",
X"b5",
X"58",
X"48",
X"10",
X"02",
X"c8",
X"c8",
X"18",
X"79",
X"d0",
X"c9",
X"95",
X"58",
X"20",
X"02",
X"bf",
X"68",
X"95",
X"58",
X"60",
X"bd",
X"96",
X"07",
X"d0",
X"1e",
X"95",
X"1e",
X"a5",
X"09",
X"29",
X"01",
X"a8",
X"c8",
X"94",
X"46",
X"88",
X"ad",
X"6a",
X"07",
X"f0",
X"02",
X"c8",
X"c8",
X"b9",
X"d4",
X"c9",
X"95",
X"58",
X"60",
X"20",
X"63",
X"bf",
X"4c",
X"02",
X"bf",
X"c9",
X"0e",
X"d0",
X"09",
X"b5",
X"16",
X"c9",
X"06",
X"d0",
X"03",
X"20",
X"98",
X"c9",
X"60",
X"20",
X"92",
X"bf",
X"4c",
X"02",
X"bf",
X"b5",
X"a0",
X"1d",
X"34",
X"04",
X"d0",
X"13",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"dd",
X"01",
X"04",
X"b0",
X"09",
X"a5",
X"09",
X"29",
X"07",
X"d0",
X"02",
X"f6",
X"cf",
X"60",
X"b5",
X"cf",
X"d5",
X"58",
X"90",
X"03",
X"4c",
X"75",
X"bf",
X"4c",
X"70",
X"bf",
X"20",
X"45",
X"cb",
X"20",
X"66",
X"cb",
X"a0",
X"01",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"11",
X"a5",
X"09",
X"29",
X"40",
X"d0",
X"02",
X"a0",
X"ff",
X"84",
X"00",
X"b5",
X"cf",
X"18",
X"65",
X"00",
X"95",
X"cf",
X"60",
X"a9",
X"13",
X"85",
X"01",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"0d",
X"b4",
X"58",
X"b5",
X"a0",
X"4a",
X"b0",
X"0a",
X"c4",
X"01",
X"f0",
X"03",
X"f6",
X"58",
X"60",
X"f6",
X"a0",
X"60",
X"98",
X"f0",
X"fa",
X"d6",
X"58",
X"60",
X"b5",
X"58",
X"48",
X"a0",
X"01",
X"b5",
X"a0",
X"29",
X"02",
X"d0",
X"0b",
X"b5",
X"58",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"95",
X"58",
X"a0",
X"02",
X"94",
X"46",
X"20",
X"02",
X"bf",
X"85",
X"00",
X"68",
X"95",
X"58",
X"60",
X"3f",
X"03",
X"b5",
X"1e",
X"29",
X"20",
X"d0",
X"4d",
X"ac",
X"cc",
X"06",
X"bd",
X"a8",
X"07",
X"39",
X"87",
X"cb",
X"d0",
X"12",
X"8a",
X"4a",
X"90",
X"04",
X"a4",
X"45",
X"b0",
X"08",
X"a0",
X"02",
X"20",
X"43",
X"e1",
X"10",
X"01",
X"88",
X"94",
X"46",
X"20",
X"df",
X"cb",
X"b5",
X"cf",
X"38",
X"fd",
X"34",
X"04",
X"c9",
X"20",
X"90",
X"02",
X"95",
X"cf",
X"b4",
X"46",
X"88",
X"d0",
X"0e",
X"b5",
X"87",
X"18",
X"75",
X"58",
X"95",
X"87",
X"b5",
X"6e",
X"69",
X"00",
X"95",
X"6e",
X"60",
X"b5",
X"87",
X"38",
X"f5",
X"58",
X"95",
X"87",
X"b5",
X"6e",
X"e9",
X"00",
X"95",
X"6e",
X"60",
X"4c",
X"8c",
X"bf",
X"b5",
X"a0",
X"29",
X"02",
X"d0",
X"37",
X"a5",
X"09",
X"29",
X"07",
X"48",
X"b5",
X"a0",
X"4a",
X"b0",
X"15",
X"68",
X"d0",
X"11",
X"bd",
X"34",
X"04",
X"18",
X"69",
X"01",
X"9d",
X"34",
X"04",
X"95",
X"58",
X"c9",
X"02",
X"d0",
X"02",
X"f6",
X"a0",
X"60",
X"68",
X"d0",
X"14",
X"bd",
X"34",
X"04",
X"38",
X"e9",
X"01",
X"9d",
X"34",
X"04",
X"95",
X"58",
X"d0",
X"07",
X"f6",
X"a0",
X"a9",
X"02",
X"9d",
X"96",
X"07",
X"60",
X"bd",
X"96",
X"07",
X"f0",
X"08",
X"a5",
X"09",
X"4a",
X"b0",
X"02",
X"f6",
X"cf",
X"60",
X"b5",
X"cf",
X"69",
X"10",
X"c5",
X"ce",
X"90",
X"f0",
X"a9",
X"00",
X"95",
X"a0",
X"60",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"03",
X"4c",
X"92",
X"bf",
X"a9",
X"e8",
X"95",
X"58",
X"4c",
X"02",
X"bf",
X"40",
X"80",
X"04",
X"04",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"03",
X"4c",
X"8c",
X"bf",
X"85",
X"03",
X"b5",
X"16",
X"38",
X"e9",
X"0a",
X"a8",
X"b9",
X"46",
X"cc",
X"85",
X"02",
X"bd",
X"01",
X"04",
X"38",
X"e5",
X"02",
X"9d",
X"01",
X"04",
X"b5",
X"87",
X"e9",
X"00",
X"95",
X"87",
X"b5",
X"6e",
X"e9",
X"00",
X"95",
X"6e",
X"a9",
X"20",
X"85",
X"02",
X"e0",
X"02",
X"90",
X"49",
X"b5",
X"58",
X"c9",
X"10",
X"90",
X"16",
X"bd",
X"17",
X"04",
X"18",
X"65",
X"02",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"65",
X"03",
X"95",
X"cf",
X"b5",
X"b6",
X"69",
X"00",
X"4c",
X"ac",
X"cc",
X"bd",
X"17",
X"04",
X"38",
X"e5",
X"02",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"e5",
X"03",
X"95",
X"cf",
X"b5",
X"b6",
X"e9",
X"00",
X"95",
X"b6",
X"a0",
X"00",
X"b5",
X"cf",
X"38",
X"fd",
X"34",
X"04",
X"10",
X"07",
X"a0",
X"10",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"c9",
X"0f",
X"90",
X"03",
X"98",
X"95",
X"58",
X"60",
X"00",
X"01",
X"03",
X"04",
X"05",
X"06",
X"07",
X"07",
X"08",
X"00",
X"03",
X"06",
X"09",
X"0b",
X"0d",
X"0e",
X"0f",
X"10",
X"00",
X"04",
X"09",
X"0d",
X"10",
X"13",
X"16",
X"17",
X"18",
X"00",
X"06",
X"0c",
X"12",
X"16",
X"1a",
X"1d",
X"1f",
X"20",
X"00",
X"07",
X"0f",
X"16",
X"1c",
X"21",
X"25",
X"27",
X"28",
X"00",
X"09",
X"12",
X"1b",
X"21",
X"27",
X"2c",
X"2f",
X"30",
X"00",
X"0b",
X"15",
X"1f",
X"27",
X"2e",
X"33",
X"37",
X"38",
X"00",
X"0c",
X"18",
X"24",
X"2d",
X"35",
X"3b",
X"3e",
X"40",
X"00",
X"0e",
X"1b",
X"28",
X"32",
X"3b",
X"42",
X"46",
X"48",
X"00",
X"0f",
X"1f",
X"2d",
X"38",
X"42",
X"4a",
X"4e",
X"50",
X"00",
X"11",
X"22",
X"31",
X"3e",
X"49",
X"51",
X"56",
X"58",
X"01",
X"03",
X"02",
X"00",
X"00",
X"09",
X"12",
X"1b",
X"24",
X"2d",
X"36",
X"3f",
X"48",
X"51",
X"5a",
X"63",
X"0c",
X"18",
X"20",
X"af",
X"f1",
X"ad",
X"d1",
X"03",
X"29",
X"08",
X"d0",
X"74",
X"ad",
X"47",
X"07",
X"d0",
X"0a",
X"bd",
X"88",
X"03",
X"20",
X"10",
X"d4",
X"29",
X"1f",
X"95",
X"a0",
X"b5",
X"a0",
X"b4",
X"16",
X"c0",
X"1f",
X"90",
X"0d",
X"c9",
X"08",
X"f0",
X"04",
X"c9",
X"18",
X"d0",
X"05",
X"18",
X"69",
X"01",
X"95",
X"a0",
X"85",
X"ef",
X"20",
X"52",
X"f1",
X"20",
X"8e",
X"ce",
X"bc",
X"e5",
X"06",
X"ad",
X"b9",
X"03",
X"99",
X"00",
X"02",
X"85",
X"07",
X"ad",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"85",
X"06",
X"a9",
X"01",
X"85",
X"00",
X"20",
X"08",
X"ce",
X"a0",
X"05",
X"b5",
X"16",
X"c9",
X"1f",
X"90",
X"02",
X"a0",
X"0b",
X"84",
X"ed",
X"a9",
X"00",
X"85",
X"00",
X"a5",
X"ef",
X"20",
X"8e",
X"ce",
X"20",
X"bb",
X"cd",
X"a5",
X"00",
X"c9",
X"04",
X"d0",
X"08",
X"ac",
X"cf",
X"06",
X"b9",
X"e5",
X"06",
X"85",
X"06",
X"e6",
X"00",
X"a5",
X"00",
X"c5",
X"ed",
X"90",
X"e2",
X"60",
X"a5",
X"03",
X"85",
X"05",
X"a4",
X"06",
X"a5",
X"01",
X"46",
X"05",
X"b0",
X"04",
X"49",
X"ff",
X"69",
X"01",
X"18",
X"6d",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"85",
X"06",
X"cd",
X"ae",
X"03",
X"b0",
X"09",
X"ad",
X"ae",
X"03",
X"38",
X"e5",
X"06",
X"4c",
X"e6",
X"cd",
X"38",
X"ed",
X"ae",
X"03",
X"c9",
X"59",
X"90",
X"04",
X"a9",
X"f8",
X"d0",
X"15",
X"ad",
X"b9",
X"03",
X"c9",
X"f8",
X"f0",
X"0e",
X"a5",
X"02",
X"46",
X"05",
X"b0",
X"04",
X"49",
X"ff",
X"69",
X"01",
X"18",
X"6d",
X"b9",
X"03",
X"99",
X"00",
X"02",
X"85",
X"07",
X"20",
X"ed",
X"ec",
X"98",
X"48",
X"ad",
X"9f",
X"07",
X"0d",
X"47",
X"07",
X"d0",
X"70",
X"85",
X"05",
X"a4",
X"b5",
X"88",
X"d0",
X"69",
X"a4",
X"ce",
X"ad",
X"54",
X"07",
X"d0",
X"05",
X"ad",
X"14",
X"07",
X"f0",
X"09",
X"e6",
X"05",
X"e6",
X"05",
X"98",
X"18",
X"69",
X"18",
X"a8",
X"98",
X"38",
X"e5",
X"07",
X"10",
X"05",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"c9",
X"08",
X"b0",
X"1c",
X"a5",
X"06",
X"c9",
X"f0",
X"b0",
X"16",
X"ad",
X"07",
X"02",
X"18",
X"69",
X"04",
X"85",
X"04",
X"38",
X"e5",
X"06",
X"10",
X"05",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"c9",
X"08",
X"90",
X"13",
X"a5",
X"05",
X"c9",
X"02",
X"f0",
X"23",
X"a4",
X"05",
X"a5",
X"ce",
X"18",
X"79",
X"3a",
X"cd",
X"e6",
X"05",
X"4c",
X"32",
X"ce",
X"a2",
X"01",
X"a5",
X"04",
X"c5",
X"06",
X"b0",
X"01",
X"e8",
X"86",
X"46",
X"a2",
X"00",
X"a5",
X"00",
X"48",
X"20",
X"2c",
X"d9",
X"68",
X"85",
X"00",
X"68",
X"18",
X"69",
X"04",
X"85",
X"06",
X"a6",
X"08",
X"60",
X"48",
X"29",
X"0f",
X"c9",
X"09",
X"90",
X"05",
X"49",
X"0f",
X"18",
X"69",
X"01",
X"85",
X"01",
X"a4",
X"00",
X"b9",
X"2e",
X"cd",
X"18",
X"65",
X"01",
X"a8",
X"b9",
X"c7",
X"cc",
X"85",
X"01",
X"68",
X"48",
X"18",
X"69",
X"08",
X"29",
X"0f",
X"c9",
X"09",
X"90",
X"05",
X"49",
X"0f",
X"18",
X"69",
X"01",
X"85",
X"02",
X"a4",
X"00",
X"b9",
X"2e",
X"cd",
X"18",
X"65",
X"02",
X"a8",
X"b9",
X"c7",
X"cc",
X"85",
X"02",
X"68",
X"4a",
X"4a",
X"4a",
X"a8",
X"b9",
X"2a",
X"cd",
X"85",
X"03",
X"60",
X"f8",
X"a0",
X"70",
X"bd",
X"00",
X"20",
X"20",
X"20",
X"00",
X"00",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"08",
X"a9",
X"00",
X"9d",
X"c5",
X"03",
X"4c",
X"92",
X"bf",
X"20",
X"02",
X"bf",
X"a0",
X"0d",
X"a9",
X"05",
X"20",
X"96",
X"bf",
X"bd",
X"34",
X"04",
X"4a",
X"4a",
X"4a",
X"4a",
X"a8",
X"b5",
X"cf",
X"38",
X"f9",
X"d5",
X"ce",
X"10",
X"05",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"c9",
X"08",
X"b0",
X"0e",
X"bd",
X"34",
X"04",
X"18",
X"69",
X"10",
X"9d",
X"34",
X"04",
X"4a",
X"4a",
X"4a",
X"4a",
X"a8",
X"b9",
X"da",
X"ce",
X"9d",
X"c5",
X"03",
X"60",
X"15",
X"30",
X"40",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"03",
X"4c",
X"63",
X"bf",
X"b5",
X"1e",
X"f0",
X"0b",
X"a9",
X"00",
X"95",
X"a0",
X"8d",
X"cb",
X"06",
X"a9",
X"10",
X"d0",
X"13",
X"a9",
X"12",
X"8d",
X"cb",
X"06",
X"a0",
X"02",
X"b9",
X"25",
X"cf",
X"99",
X"01",
X"00",
X"88",
X"10",
X"f7",
X"20",
X"6c",
X"cf",
X"95",
X"58",
X"a0",
X"01",
X"b5",
X"a0",
X"29",
X"01",
X"d0",
X"0a",
X"b5",
X"58",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"95",
X"58",
X"c8",
X"94",
X"46",
X"4c",
X"02",
X"bf",
X"a0",
X"00",
X"20",
X"43",
X"e1",
X"10",
X"0a",
X"c8",
X"a5",
X"00",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"00",
X"a5",
X"00",
X"c9",
X"3c",
X"90",
X"1c",
X"a9",
X"3c",
X"85",
X"00",
X"b5",
X"16",
X"c9",
X"11",
X"d0",
X"12",
X"98",
X"d5",
X"a0",
X"f0",
X"0d",
X"b5",
X"a0",
X"f0",
X"06",
X"d6",
X"58",
X"b5",
X"58",
X"d0",
X"40",
X"98",
X"95",
X"a0",
X"a5",
X"00",
X"29",
X"3c",
X"4a",
X"4a",
X"85",
X"00",
X"a0",
X"00",
X"a5",
X"57",
X"f0",
X"24",
X"ad",
X"75",
X"07",
X"f0",
X"1f",
X"c8",
X"a5",
X"57",
X"c9",
X"19",
X"90",
X"08",
X"ad",
X"75",
X"07",
X"c9",
X"02",
X"90",
X"01",
X"c8",
X"b5",
X"16",
X"c9",
X"12",
X"d0",
X"04",
X"a5",
X"57",
X"d0",
X"06",
X"b5",
X"a0",
X"d0",
X"02",
X"a0",
X"00",
X"b9",
X"01",
X"00",
X"a4",
X"00",
X"38",
X"e9",
X"01",
X"88",
X"10",
X"fa",
X"60",
X"1a",
X"58",
X"98",
X"96",
X"94",
X"92",
X"90",
X"8e",
X"8c",
X"8a",
X"88",
X"86",
X"84",
X"82",
X"80",
X"ae",
X"68",
X"03",
X"b5",
X"16",
X"c9",
X"2d",
X"d0",
X"10",
X"86",
X"08",
X"b5",
X"1e",
X"f0",
X"1a",
X"29",
X"40",
X"f0",
X"06",
X"b5",
X"cf",
X"c9",
X"e0",
X"90",
X"0a",
X"a9",
X"80",
X"85",
X"fc",
X"ee",
X"72",
X"07",
X"4c",
X"71",
X"d0",
X"20",
X"8c",
X"bf",
X"4c",
X"7b",
X"d1",
X"ce",
X"64",
X"03",
X"d0",
X"44",
X"a9",
X"04",
X"8d",
X"64",
X"03",
X"ad",
X"63",
X"03",
X"49",
X"01",
X"8d",
X"63",
X"03",
X"a9",
X"22",
X"85",
X"05",
X"ac",
X"69",
X"03",
X"b9",
X"dd",
X"cf",
X"85",
X"04",
X"ac",
X"00",
X"03",
X"c8",
X"a2",
X"0c",
X"20",
X"cd",
X"8a",
X"a6",
X"08",
X"20",
X"8f",
X"8a",
X"a9",
X"08",
X"85",
X"fe",
X"a9",
X"01",
X"85",
X"fd",
X"ee",
X"69",
X"03",
X"ad",
X"69",
X"03",
X"c9",
X"0f",
X"d0",
X"0b",
X"20",
X"63",
X"c3",
X"a9",
X"40",
X"95",
X"1e",
X"a9",
X"80",
X"85",
X"fe",
X"4c",
X"7b",
X"d1",
X"21",
X"41",
X"11",
X"31",
X"b5",
X"1e",
X"29",
X"20",
X"f0",
X"14",
X"b5",
X"cf",
X"c9",
X"e0",
X"90",
X"9e",
X"a2",
X"04",
X"20",
X"98",
X"c9",
X"ca",
X"10",
X"fa",
X"8d",
X"cb",
X"06",
X"a6",
X"08",
X"60",
X"a9",
X"00",
X"8d",
X"cb",
X"06",
X"ad",
X"47",
X"07",
X"f0",
X"03",
X"4c",
X"39",
X"d1",
X"ad",
X"63",
X"03",
X"10",
X"03",
X"4c",
X"0f",
X"d1",
X"ce",
X"64",
X"03",
X"d0",
X"0d",
X"a9",
X"20",
X"8d",
X"64",
X"03",
X"ad",
X"63",
X"03",
X"49",
X"01",
X"8d",
X"63",
X"03",
X"a5",
X"09",
X"29",
X"0f",
X"d0",
X"04",
X"a9",
X"02",
X"95",
X"46",
X"bd",
X"8a",
X"07",
X"f0",
X"1c",
X"20",
X"43",
X"e1",
X"10",
X"17",
X"a9",
X"01",
X"95",
X"46",
X"a9",
X"02",
X"8d",
X"65",
X"03",
X"a9",
X"20",
X"9d",
X"8a",
X"07",
X"8d",
X"90",
X"07",
X"b5",
X"87",
X"c9",
X"c8",
X"b0",
X"3e",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"38",
X"b5",
X"87",
X"cd",
X"66",
X"03",
X"d0",
X"0c",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"a8",
X"b9",
X"61",
X"d0",
X"8d",
X"dc",
X"06",
X"b5",
X"87",
X"18",
X"6d",
X"65",
X"03",
X"95",
X"87",
X"b4",
X"46",
X"c0",
X"01",
X"f0",
X"17",
X"a0",
X"ff",
X"38",
X"ed",
X"66",
X"03",
X"10",
X"07",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"a0",
X"01",
X"cd",
X"dc",
X"06",
X"90",
X"03",
X"8c",
X"65",
X"03",
X"bd",
X"8a",
X"07",
X"d0",
X"28",
X"20",
X"8c",
X"bf",
X"ad",
X"5f",
X"07",
X"c9",
X"05",
X"90",
X"09",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"03",
X"20",
X"94",
X"ba",
X"b5",
X"cf",
X"c9",
X"80",
X"90",
X"1c",
X"bd",
X"a7",
X"07",
X"29",
X"03",
X"a8",
X"b9",
X"61",
X"d0",
X"9d",
X"8a",
X"07",
X"4c",
X"49",
X"d1",
X"c9",
X"01",
X"d0",
X"09",
X"d6",
X"cf",
X"20",
X"63",
X"c3",
X"a9",
X"fe",
X"95",
X"a0",
X"ad",
X"5f",
X"07",
X"c9",
X"07",
X"f0",
X"04",
X"c9",
X"05",
X"b0",
X"27",
X"ad",
X"90",
X"07",
X"d0",
X"22",
X"a9",
X"20",
X"8d",
X"90",
X"07",
X"ad",
X"63",
X"03",
X"49",
X"80",
X"8d",
X"63",
X"03",
X"30",
X"e1",
X"20",
X"d9",
X"d1",
X"ac",
X"cc",
X"06",
X"f0",
X"03",
X"38",
X"e9",
X"10",
X"8d",
X"90",
X"07",
X"a9",
X"15",
X"8d",
X"cb",
X"06",
X"20",
X"bc",
X"d1",
X"a0",
X"10",
X"b5",
X"46",
X"4a",
X"90",
X"02",
X"a0",
X"f0",
X"98",
X"18",
X"75",
X"87",
X"ac",
X"cf",
X"06",
X"99",
X"87",
X"00",
X"b5",
X"cf",
X"18",
X"69",
X"08",
X"99",
X"cf",
X"00",
X"b5",
X"1e",
X"99",
X"1e",
X"00",
X"b5",
X"46",
X"99",
X"46",
X"00",
X"a5",
X"08",
X"48",
X"ae",
X"cf",
X"06",
X"86",
X"08",
X"a9",
X"2d",
X"95",
X"16",
X"20",
X"bc",
X"d1",
X"68",
X"85",
X"08",
X"aa",
X"a9",
X"00",
X"8d",
X"6a",
X"03",
X"60",
X"ee",
X"6a",
X"03",
X"20",
X"d7",
X"c8",
X"b5",
X"1e",
X"d0",
X"f5",
X"a9",
X"0a",
X"9d",
X"9a",
X"04",
X"20",
X"43",
X"e2",
X"4c",
X"53",
X"d8",
X"bf",
X"40",
X"bf",
X"bf",
X"bf",
X"40",
X"40",
X"bf",
X"ac",
X"67",
X"03",
X"ee",
X"67",
X"03",
X"ad",
X"67",
X"03",
X"29",
X"07",
X"8d",
X"67",
X"03",
X"b9",
X"d1",
X"d1",
X"60",
X"ad",
X"47",
X"07",
X"d0",
X"30",
X"a9",
X"40",
X"ac",
X"cc",
X"06",
X"f0",
X"02",
X"a9",
X"60",
X"85",
X"00",
X"bd",
X"01",
X"04",
X"38",
X"e5",
X"00",
X"9d",
X"01",
X"04",
X"b5",
X"87",
X"e9",
X"01",
X"95",
X"87",
X"b5",
X"6e",
X"e9",
X"00",
X"95",
X"6e",
X"bc",
X"17",
X"04",
X"b5",
X"cf",
X"d9",
X"9d",
X"c5",
X"f0",
X"06",
X"18",
X"7d",
X"34",
X"04",
X"95",
X"cf",
X"20",
X"52",
X"f1",
X"b5",
X"1e",
X"d0",
X"c3",
X"a9",
X"51",
X"85",
X"00",
X"a0",
X"02",
X"a5",
X"09",
X"29",
X"02",
X"f0",
X"02",
X"a0",
X"82",
X"84",
X"01",
X"bc",
X"e5",
X"06",
X"a2",
X"00",
X"ad",
X"b9",
X"03",
X"99",
X"00",
X"02",
X"a5",
X"00",
X"99",
X"01",
X"02",
X"e6",
X"00",
X"a5",
X"01",
X"99",
X"02",
X"02",
X"ad",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"18",
X"69",
X"08",
X"8d",
X"ae",
X"03",
X"c8",
X"c8",
X"c8",
X"c8",
X"e8",
X"e0",
X"03",
X"90",
X"d9",
X"a6",
X"08",
X"20",
X"af",
X"f1",
X"bc",
X"e5",
X"06",
X"ad",
X"d1",
X"03",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"0c",
X"02",
X"68",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"08",
X"02",
X"68",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"04",
X"02",
X"68",
X"4a",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"60",
X"d6",
X"a0",
X"d0",
X"0c",
X"a9",
X"08",
X"95",
X"a0",
X"f6",
X"58",
X"b5",
X"58",
X"c9",
X"03",
X"b0",
X"18",
X"20",
X"52",
X"f1",
X"ad",
X"b9",
X"03",
X"8d",
X"ba",
X"03",
X"ad",
X"ae",
X"03",
X"8d",
X"af",
X"03",
X"bc",
X"e5",
X"06",
X"b5",
X"58",
X"20",
X"17",
X"ed",
X"60",
X"a9",
X"00",
X"95",
X"0f",
X"a9",
X"08",
X"85",
X"fe",
X"a9",
X"05",
X"8d",
X"38",
X"01",
X"4c",
X"36",
X"d3",
X"00",
X"00",
X"08",
X"08",
X"00",
X"08",
X"00",
X"08",
X"54",
X"55",
X"56",
X"57",
X"a9",
X"00",
X"8d",
X"cb",
X"06",
X"ad",
X"46",
X"07",
X"c9",
X"05",
X"b0",
X"2c",
X"20",
X"04",
X"8e",
X"11",
X"d3",
X"f2",
X"d2",
X"12",
X"d3",
X"4e",
X"d3",
X"a2",
X"d3",
X"a0",
X"05",
X"ad",
X"fa",
X"07",
X"c9",
X"01",
X"f0",
X"0e",
X"a0",
X"03",
X"c9",
X"03",
X"f0",
X"08",
X"a0",
X"00",
X"c9",
X"06",
X"f0",
X"02",
X"a9",
X"ff",
X"8d",
X"d7",
X"06",
X"94",
X"1e",
X"ee",
X"46",
X"07",
X"60",
X"ad",
X"f8",
X"07",
X"0d",
X"f9",
X"07",
X"0d",
X"fa",
X"07",
X"f0",
X"f1",
X"a5",
X"09",
X"29",
X"04",
X"f0",
X"04",
X"a9",
X"10",
X"85",
X"fe",
X"a0",
X"23",
X"a9",
X"ff",
X"8d",
X"39",
X"01",
X"20",
X"5f",
X"8f",
X"a9",
X"05",
X"8d",
X"39",
X"01",
X"a0",
X"0b",
X"ad",
X"53",
X"07",
X"f0",
X"02",
X"a0",
X"11",
X"20",
X"5f",
X"8f",
X"ad",
X"53",
X"07",
X"0a",
X"0a",
X"0a",
X"0a",
X"09",
X"04",
X"4c",
X"36",
X"bc",
X"b5",
X"cf",
X"c9",
X"72",
X"90",
X"05",
X"d6",
X"cf",
X"4c",
X"65",
X"d3",
X"ad",
X"d7",
X"06",
X"f0",
X"38",
X"30",
X"36",
X"a9",
X"16",
X"8d",
X"cb",
X"06",
X"20",
X"52",
X"f1",
X"bc",
X"e5",
X"06",
X"a2",
X"03",
X"ad",
X"b9",
X"03",
X"18",
X"7d",
X"cd",
X"d2",
X"99",
X"00",
X"02",
X"bd",
X"d5",
X"d2",
X"99",
X"01",
X"02",
X"a9",
X"22",
X"99",
X"02",
X"02",
X"ad",
X"ae",
X"03",
X"18",
X"7d",
X"d1",
X"d2",
X"99",
X"03",
X"02",
X"c8",
X"c8",
X"c8",
X"c8",
X"ca",
X"10",
X"da",
X"a6",
X"08",
X"60",
X"20",
X"65",
X"d3",
X"a9",
X"06",
X"9d",
X"96",
X"07",
X"ee",
X"46",
X"07",
X"60",
X"20",
X"65",
X"d3",
X"bd",
X"96",
X"07",
X"d0",
X"05",
X"ad",
X"b1",
X"07",
X"f0",
X"ef",
X"60",
X"b5",
X"1e",
X"d0",
X"56",
X"bd",
X"8a",
X"07",
X"d0",
X"51",
X"b5",
X"a0",
X"d0",
X"23",
X"b5",
X"58",
X"30",
X"14",
X"20",
X"43",
X"e1",
X"10",
X"09",
X"a5",
X"00",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"85",
X"00",
X"a5",
X"00",
X"c9",
X"21",
X"90",
X"35",
X"b5",
X"58",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"95",
X"58",
X"f6",
X"a0",
X"bd",
X"34",
X"04",
X"b4",
X"58",
X"10",
X"03",
X"bd",
X"17",
X"04",
X"85",
X"00",
X"a5",
X"09",
X"4a",
X"90",
X"19",
X"ad",
X"47",
X"07",
X"d0",
X"14",
X"b5",
X"cf",
X"18",
X"75",
X"58",
X"95",
X"cf",
X"c5",
X"00",
X"d0",
X"09",
X"a9",
X"00",
X"95",
X"a0",
X"a9",
X"40",
X"9d",
X"8a",
X"07",
X"a9",
X"20",
X"9d",
X"c5",
X"03",
X"60",
X"85",
X"07",
X"b5",
X"34",
X"d0",
X"0e",
X"a0",
X"18",
X"b5",
X"58",
X"18",
X"65",
X"07",
X"95",
X"58",
X"b5",
X"a0",
X"69",
X"00",
X"60",
X"a0",
X"08",
X"b5",
X"58",
X"38",
X"e5",
X"07",
X"95",
X"58",
X"b5",
X"a0",
X"e9",
X"00",
X"60",
X"b5",
X"b6",
X"c9",
X"03",
X"d0",
X"03",
X"4c",
X"98",
X"c9",
X"b5",
X"1e",
X"10",
X"01",
X"60",
X"a8",
X"bd",
X"a2",
X"03",
X"85",
X"00",
X"b5",
X"46",
X"f0",
X"03",
X"4c",
X"bb",
X"d5",
X"a9",
X"2d",
X"d5",
X"cf",
X"90",
X"0f",
X"c4",
X"00",
X"f0",
X"08",
X"18",
X"69",
X"02",
X"95",
X"cf",
X"4c",
X"b1",
X"d5",
X"4c",
X"98",
X"d5",
X"d9",
X"cf",
X"00",
X"90",
X"0d",
X"e4",
X"00",
X"f0",
X"f4",
X"18",
X"69",
X"02",
X"99",
X"cf",
X"00",
X"4c",
X"b1",
X"d5",
X"b5",
X"cf",
X"48",
X"bd",
X"a2",
X"03",
X"10",
X"18",
X"bd",
X"34",
X"04",
X"18",
X"69",
X"05",
X"85",
X"00",
X"b5",
X"a0",
X"69",
X"00",
X"30",
X"1a",
X"d0",
X"0c",
X"a5",
X"00",
X"c9",
X"0b",
X"90",
X"0c",
X"b0",
X"04",
X"c5",
X"08",
X"f0",
X"0c",
X"20",
X"b7",
X"bf",
X"4c",
X"a7",
X"d4",
X"20",
X"b1",
X"d5",
X"4c",
X"a7",
X"d4",
X"20",
X"b4",
X"bf",
X"b4",
X"1e",
X"68",
X"38",
X"f5",
X"cf",
X"18",
X"79",
X"cf",
X"00",
X"99",
X"cf",
X"00",
X"bd",
X"a2",
X"03",
X"30",
X"04",
X"aa",
X"20",
X"21",
X"dc",
X"a4",
X"08",
X"b9",
X"a0",
X"00",
X"19",
X"34",
X"04",
X"f0",
X"77",
X"ae",
X"00",
X"03",
X"e0",
X"20",
X"b0",
X"70",
X"b9",
X"a0",
X"00",
X"48",
X"48",
X"20",
X"41",
X"d5",
X"a5",
X"01",
X"9d",
X"01",
X"03",
X"a5",
X"00",
X"9d",
X"02",
X"03",
X"a9",
X"02",
X"9d",
X"03",
X"03",
X"b9",
X"a0",
X"00",
X"30",
X"0d",
X"a9",
X"a2",
X"9d",
X"04",
X"03",
X"a9",
X"a3",
X"9d",
X"05",
X"03",
X"4c",
X"ff",
X"d4",
X"a9",
X"24",
X"9d",
X"04",
X"03",
X"9d",
X"05",
X"03",
X"b9",
X"1e",
X"00",
X"a8",
X"68",
X"49",
X"ff",
X"20",
X"41",
X"d5",
X"a5",
X"01",
X"9d",
X"06",
X"03",
X"a5",
X"00",
X"9d",
X"07",
X"03",
X"a9",
X"02",
X"9d",
X"08",
X"03",
X"68",
X"10",
X"0d",
X"a9",
X"a2",
X"9d",
X"09",
X"03",
X"a9",
X"a3",
X"9d",
X"0a",
X"03",
X"4c",
X"30",
X"d5",
X"a9",
X"24",
X"9d",
X"09",
X"03",
X"9d",
X"0a",
X"03",
X"a9",
X"00",
X"9d",
X"0b",
X"03",
X"ad",
X"00",
X"03",
X"18",
X"69",
X"0a",
X"8d",
X"00",
X"03",
X"a6",
X"08",
X"60",
X"48",
X"b9",
X"87",
X"00",
X"18",
X"69",
X"08",
X"ae",
X"cc",
X"06",
X"d0",
X"03",
X"18",
X"69",
X"10",
X"48",
X"b9",
X"6e",
X"00",
X"69",
X"00",
X"85",
X"02",
X"68",
X"29",
X"f0",
X"4a",
X"4a",
X"4a",
X"85",
X"00",
X"b6",
X"cf",
X"68",
X"10",
X"05",
X"8a",
X"18",
X"69",
X"08",
X"aa",
X"8a",
X"ae",
X"00",
X"03",
X"0a",
X"2a",
X"48",
X"2a",
X"29",
X"03",
X"09",
X"20",
X"85",
X"01",
X"a5",
X"02",
X"29",
X"01",
X"0a",
X"0a",
X"05",
X"01",
X"85",
X"01",
X"68",
X"29",
X"e0",
X"18",
X"65",
X"00",
X"85",
X"00",
X"b9",
X"cf",
X"00",
X"c9",
X"e8",
X"90",
X"06",
X"a5",
X"00",
X"29",
X"bf",
X"85",
X"00",
X"60",
X"98",
X"aa",
X"20",
X"af",
X"f1",
X"a9",
X"06",
X"20",
X"11",
X"da",
X"ad",
X"ad",
X"03",
X"9d",
X"17",
X"01",
X"a5",
X"ce",
X"9d",
X"1e",
X"01",
X"a9",
X"01",
X"95",
X"46",
X"20",
X"63",
X"c3",
X"99",
X"a0",
X"00",
X"99",
X"34",
X"04",
X"60",
X"98",
X"48",
X"20",
X"6b",
X"bf",
X"68",
X"aa",
X"20",
X"6b",
X"bf",
X"a6",
X"08",
X"bd",
X"a2",
X"03",
X"30",
X"04",
X"aa",
X"20",
X"21",
X"dc",
X"a6",
X"08",
X"60",
X"b5",
X"a0",
X"1d",
X"34",
X"04",
X"d0",
X"15",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"dd",
X"01",
X"04",
X"b0",
X"0b",
X"a5",
X"09",
X"29",
X"07",
X"d0",
X"02",
X"f6",
X"cf",
X"4c",
X"fe",
X"d5",
X"b5",
X"cf",
X"d5",
X"58",
X"90",
X"06",
X"20",
X"b7",
X"bf",
X"4c",
X"fe",
X"d5",
X"20",
X"b4",
X"bf",
X"bd",
X"a2",
X"03",
X"30",
X"03",
X"20",
X"21",
X"dc",
X"60",
X"a9",
X"0e",
X"20",
X"47",
X"cb",
X"20",
X"66",
X"cb",
X"bd",
X"a2",
X"03",
X"30",
X"1c",
X"a5",
X"86",
X"18",
X"65",
X"00",
X"85",
X"86",
X"a5",
X"6d",
X"a4",
X"00",
X"30",
X"05",
X"69",
X"00",
X"4c",
X"28",
X"d6",
X"e9",
X"00",
X"85",
X"6d",
X"8c",
X"a1",
X"03",
X"20",
X"21",
X"dc",
X"60",
X"bd",
X"a2",
X"03",
X"30",
X"06",
X"20",
X"88",
X"bf",
X"20",
X"21",
X"dc",
X"60",
X"20",
X"02",
X"bf",
X"85",
X"00",
X"bd",
X"a2",
X"03",
X"30",
X"07",
X"a9",
X"10",
X"95",
X"58",
X"20",
X"14",
X"d6",
X"60",
X"20",
X"5b",
X"d6",
X"4c",
X"fe",
X"d5",
X"20",
X"5b",
X"d6",
X"4c",
X"71",
X"d6",
X"ad",
X"47",
X"07",
X"d0",
X"19",
X"bd",
X"17",
X"04",
X"18",
X"7d",
X"34",
X"04",
X"9d",
X"17",
X"04",
X"b5",
X"cf",
X"75",
X"a0",
X"95",
X"cf",
X"60",
X"bd",
X"a2",
X"03",
X"f0",
X"03",
X"20",
X"19",
X"dc",
X"60",
X"b5",
X"16",
X"c9",
X"14",
X"f0",
X"55",
X"ad",
X"1c",
X"07",
X"b4",
X"16",
X"c0",
X"05",
X"f0",
X"04",
X"c0",
X"0d",
X"d0",
X"02",
X"69",
X"38",
X"e9",
X"48",
X"85",
X"01",
X"ad",
X"1a",
X"07",
X"e9",
X"00",
X"85",
X"00",
X"ad",
X"1d",
X"07",
X"69",
X"48",
X"85",
X"03",
X"ad",
X"1b",
X"07",
X"69",
X"00",
X"85",
X"02",
X"b5",
X"87",
X"c5",
X"01",
X"b5",
X"6e",
X"e5",
X"00",
X"30",
X"20",
X"b5",
X"87",
X"c5",
X"03",
X"b5",
X"6e",
X"e5",
X"02",
X"30",
X"19",
X"b5",
X"1e",
X"c9",
X"05",
X"f0",
X"13",
X"c0",
X"0d",
X"f0",
X"0f",
X"c0",
X"30",
X"f0",
X"0b",
X"c0",
X"31",
X"f0",
X"07",
X"c0",
X"32",
X"f0",
X"03",
X"20",
X"98",
X"c9",
X"60",
X"ff",
X"ff",
X"ff",
X"b5",
X"24",
X"f0",
X"56",
X"0a",
X"b0",
X"53",
X"a5",
X"09",
X"4a",
X"b0",
X"4e",
X"8a",
X"0a",
X"0a",
X"18",
X"69",
X"1c",
X"a8",
X"a2",
X"04",
X"86",
X"01",
X"98",
X"48",
X"b5",
X"1e",
X"29",
X"20",
X"d0",
X"34",
X"b5",
X"0f",
X"f0",
X"30",
X"b5",
X"16",
X"c9",
X"24",
X"90",
X"04",
X"c9",
X"2b",
X"90",
X"26",
X"c9",
X"06",
X"d0",
X"06",
X"b5",
X"1e",
X"c9",
X"02",
X"b0",
X"1c",
X"bd",
X"d8",
X"03",
X"d0",
X"17",
X"8a",
X"0a",
X"0a",
X"18",
X"69",
X"04",
X"aa",
X"20",
X"27",
X"e3",
X"a6",
X"08",
X"90",
X"09",
X"a9",
X"80",
X"95",
X"24",
X"a6",
X"01",
X"20",
X"3e",
X"d7",
X"68",
X"a8",
X"a6",
X"01",
X"ca",
X"10",
X"bb",
X"a6",
X"08",
X"60",
X"06",
X"00",
X"02",
X"12",
X"11",
X"07",
X"05",
X"2d",
X"20",
X"52",
X"f1",
X"a6",
X"01",
X"b5",
X"0f",
X"10",
X"0b",
X"29",
X"0f",
X"aa",
X"b5",
X"16",
X"c9",
X"2d",
X"f0",
X"0c",
X"a6",
X"01",
X"b5",
X"16",
X"c9",
X"02",
X"f0",
X"6b",
X"c9",
X"2d",
X"d0",
X"2d",
X"ce",
X"83",
X"04",
X"d0",
X"62",
X"20",
X"63",
X"c3",
X"95",
X"58",
X"8d",
X"cb",
X"06",
X"a9",
X"fe",
X"95",
X"a0",
X"ac",
X"5f",
X"07",
X"b9",
X"36",
X"d7",
X"95",
X"16",
X"a9",
X"20",
X"c0",
X"03",
X"b0",
X"02",
X"09",
X"03",
X"95",
X"1e",
X"a9",
X"80",
X"85",
X"fe",
X"a6",
X"01",
X"a9",
X"09",
X"d0",
X"33",
X"c9",
X"08",
X"f0",
X"36",
X"c9",
X"0c",
X"f0",
X"32",
X"c9",
X"15",
X"b0",
X"2e",
X"b5",
X"16",
X"c9",
X"0d",
X"d0",
X"06",
X"b5",
X"cf",
X"69",
X"18",
X"95",
X"cf",
X"20",
X"1b",
X"e0",
X"b5",
X"1e",
X"29",
X"1f",
X"09",
X"20",
X"95",
X"1e",
X"a9",
X"02",
X"b4",
X"16",
X"c0",
X"05",
X"d0",
X"02",
X"a9",
X"06",
X"c0",
X"06",
X"d0",
X"02",
X"a9",
X"01",
X"20",
X"11",
X"da",
X"a9",
X"08",
X"85",
X"ff",
X"60",
X"a5",
X"09",
X"4a",
X"90",
X"36",
X"ad",
X"47",
X"07",
X"0d",
X"d6",
X"03",
X"d0",
X"2e",
X"8a",
X"0a",
X"0a",
X"18",
X"69",
X"24",
X"a8",
X"20",
X"25",
X"e3",
X"a6",
X"08",
X"90",
X"1b",
X"bd",
X"be",
X"06",
X"d0",
X"1b",
X"a9",
X"01",
X"9d",
X"be",
X"06",
X"b5",
X"64",
X"49",
X"ff",
X"18",
X"69",
X"01",
X"95",
X"64",
X"ad",
X"9f",
X"07",
X"d0",
X"08",
X"4c",
X"2c",
X"d9",
X"a9",
X"00",
X"9d",
X"be",
X"06",
X"60",
X"20",
X"98",
X"c9",
X"a9",
X"06",
X"20",
X"11",
X"da",
X"a9",
X"20",
X"85",
X"fe",
X"a5",
X"39",
X"c9",
X"02",
X"90",
X"0e",
X"c9",
X"03",
X"f0",
X"24",
X"a9",
X"23",
X"8d",
X"9f",
X"07",
X"a9",
X"40",
X"85",
X"fb",
X"60",
X"ad",
X"56",
X"07",
X"f0",
X"1b",
X"c9",
X"01",
X"d0",
X"23",
X"a6",
X"08",
X"a9",
X"02",
X"8d",
X"56",
X"07",
X"20",
X"f1",
X"85",
X"a6",
X"08",
X"a9",
X"0c",
X"4c",
X"47",
X"d8",
X"a9",
X"0b",
X"9d",
X"10",
X"01",
X"60",
X"a9",
X"01",
X"8d",
X"56",
X"07",
X"a9",
X"09",
X"a0",
X"00",
X"20",
X"48",
X"d9",
X"60",
X"18",
X"e8",
X"30",
X"d0",
X"08",
X"f8",
X"a5",
X"09",
X"4a",
X"b0",
X"f4",
X"20",
X"41",
X"dc",
X"b0",
X"23",
X"bd",
X"d8",
X"03",
X"d0",
X"1e",
X"a5",
X"0e",
X"c9",
X"08",
X"d0",
X"18",
X"b5",
X"1e",
X"29",
X"20",
X"d0",
X"12",
X"20",
X"52",
X"dc",
X"20",
X"25",
X"e3",
X"a6",
X"08",
X"b0",
X"09",
X"bd",
X"91",
X"04",
X"29",
X"fe",
X"9d",
X"91",
X"04",
X"60",
X"b4",
X"16",
X"c0",
X"2e",
X"d0",
X"03",
X"4c",
X"00",
X"d8",
X"ad",
X"9f",
X"07",
X"f0",
X"06",
X"4c",
X"95",
X"d7",
X"0a",
X"06",
X"04",
X"bd",
X"91",
X"04",
X"29",
X"01",
X"1d",
X"d8",
X"03",
X"d0",
X"59",
X"a9",
X"01",
X"1d",
X"91",
X"04",
X"9d",
X"91",
X"04",
X"c0",
X"12",
X"f0",
X"4e",
X"c0",
X"0d",
X"f0",
X"7d",
X"c0",
X"0c",
X"f0",
X"79",
X"c0",
X"33",
X"f0",
X"42",
X"c0",
X"15",
X"b0",
X"71",
X"ad",
X"4e",
X"07",
X"f0",
X"6c",
X"b5",
X"1e",
X"0a",
X"b0",
X"34",
X"b5",
X"1e",
X"29",
X"07",
X"c9",
X"02",
X"90",
X"2c",
X"b5",
X"16",
X"c9",
X"06",
X"f0",
X"25",
X"a9",
X"08",
X"85",
X"ff",
X"b5",
X"1e",
X"09",
X"80",
X"95",
X"1e",
X"20",
X"05",
X"da",
X"b9",
X"4f",
X"d8",
X"95",
X"58",
X"a9",
X"03",
X"18",
X"6d",
X"84",
X"04",
X"bc",
X"96",
X"07",
X"c0",
X"03",
X"b0",
X"03",
X"b9",
X"92",
X"d8",
X"20",
X"11",
X"da",
X"60",
X"a5",
X"9f",
X"30",
X"02",
X"d0",
X"6a",
X"b5",
X"16",
X"c9",
X"07",
X"90",
X"09",
X"a5",
X"ce",
X"18",
X"69",
X"0c",
X"d5",
X"cf",
X"90",
X"5b",
X"ad",
X"91",
X"07",
X"d0",
X"56",
X"ad",
X"9e",
X"07",
X"d0",
X"3d",
X"ad",
X"ad",
X"03",
X"cd",
X"ae",
X"03",
X"90",
X"03",
X"4c",
X"f6",
X"d9",
X"b5",
X"46",
X"c9",
X"01",
X"d0",
X"03",
X"4c",
X"ff",
X"d9",
X"ad",
X"9e",
X"07",
X"d0",
X"24",
X"ae",
X"56",
X"07",
X"f0",
X"22",
X"8d",
X"56",
X"07",
X"a9",
X"08",
X"8d",
X"9e",
X"07",
X"0a",
X"85",
X"ff",
X"20",
X"f1",
X"85",
X"a9",
X"0a",
X"a0",
X"01",
X"85",
X"0e",
X"84",
X"1d",
X"a0",
X"ff",
X"8c",
X"47",
X"07",
X"c8",
X"8c",
X"75",
X"07",
X"a6",
X"08",
X"60",
X"86",
X"57",
X"e8",
X"86",
X"fc",
X"a9",
X"fc",
X"85",
X"9f",
X"a9",
X"0b",
X"d0",
X"e1",
X"02",
X"06",
X"05",
X"06",
X"b5",
X"16",
X"c9",
X"12",
X"f0",
X"bd",
X"a9",
X"04",
X"85",
X"ff",
X"b5",
X"16",
X"a0",
X"00",
X"c9",
X"14",
X"f0",
X"1b",
X"c9",
X"08",
X"f0",
X"17",
X"c9",
X"33",
X"f0",
X"13",
X"c9",
X"0c",
X"f0",
X"0f",
X"c8",
X"c9",
X"05",
X"f0",
X"0a",
X"c8",
X"c9",
X"11",
X"f0",
X"05",
X"c8",
X"c9",
X"07",
X"d0",
X"1d",
X"b9",
X"65",
X"d9",
X"20",
X"11",
X"da",
X"b5",
X"46",
X"48",
X"20",
X"2f",
X"e0",
X"68",
X"95",
X"46",
X"a9",
X"20",
X"95",
X"1e",
X"20",
X"63",
X"c3",
X"95",
X"58",
X"a9",
X"fd",
X"85",
X"9f",
X"60",
X"c9",
X"09",
X"90",
X"1d",
X"29",
X"01",
X"95",
X"16",
X"a0",
X"00",
X"94",
X"1e",
X"a9",
X"03",
X"20",
X"11",
X"da",
X"20",
X"63",
X"c3",
X"20",
X"05",
X"da",
X"b9",
X"51",
X"d8",
X"95",
X"58",
X"4c",
X"f1",
X"d9",
X"10",
X"0b",
X"a9",
X"04",
X"95",
X"1e",
X"ee",
X"84",
X"04",
X"ad",
X"84",
X"04",
X"18",
X"6d",
X"91",
X"07",
X"20",
X"11",
X"da",
X"ee",
X"91",
X"07",
X"ac",
X"6a",
X"07",
X"b9",
X"d2",
X"d9",
X"9d",
X"96",
X"07",
X"a9",
X"fc",
X"85",
X"9f",
X"60",
X"b5",
X"46",
X"c9",
X"01",
X"d0",
X"03",
X"4c",
X"2c",
X"d9",
X"20",
X"1c",
X"db",
X"4c",
X"2c",
X"d9",
X"a0",
X"01",
X"20",
X"43",
X"e1",
X"10",
X"01",
X"c8",
X"94",
X"46",
X"88",
X"60",
X"9d",
X"10",
X"01",
X"a9",
X"30",
X"9d",
X"2c",
X"01",
X"b5",
X"cf",
X"9d",
X"1e",
X"01",
X"ad",
X"ae",
X"03",
X"9d",
X"17",
X"01",
X"60",
X"80",
X"40",
X"20",
X"10",
X"08",
X"04",
X"02",
X"7f",
X"bf",
X"df",
X"ef",
X"f7",
X"fb",
X"fd",
X"a5",
X"09",
X"4a",
X"90",
X"ec",
X"ad",
X"4e",
X"07",
X"f0",
X"e7",
X"b5",
X"16",
X"c9",
X"15",
X"b0",
X"6e",
X"c9",
X"11",
X"f0",
X"6a",
X"c9",
X"0d",
X"f0",
X"66",
X"bd",
X"d8",
X"03",
X"d0",
X"61",
X"20",
X"52",
X"dc",
X"ca",
X"30",
X"5b",
X"86",
X"01",
X"98",
X"48",
X"b5",
X"0f",
X"f0",
X"4c",
X"b5",
X"16",
X"c9",
X"15",
X"b0",
X"46",
X"c9",
X"11",
X"f0",
X"42",
X"c9",
X"0d",
X"f0",
X"3e",
X"bd",
X"d8",
X"03",
X"d0",
X"39",
X"8a",
X"0a",
X"0a",
X"18",
X"69",
X"04",
X"aa",
X"20",
X"27",
X"e3",
X"a6",
X"08",
X"a4",
X"01",
X"90",
X"20",
X"b5",
X"1e",
X"19",
X"1e",
X"00",
X"29",
X"80",
X"d0",
X"11",
X"b9",
X"91",
X"04",
X"3d",
X"25",
X"da",
X"d0",
X"18",
X"b9",
X"91",
X"04",
X"1d",
X"25",
X"da",
X"99",
X"91",
X"04",
X"20",
X"b4",
X"da",
X"4c",
X"aa",
X"da",
X"b9",
X"91",
X"04",
X"3d",
X"2c",
X"da",
X"99",
X"91",
X"04",
X"68",
X"a8",
X"a6",
X"01",
X"ca",
X"10",
X"a5",
X"a6",
X"08",
X"60",
X"b9",
X"1e",
X"00",
X"15",
X"1e",
X"29",
X"20",
X"d0",
X"33",
X"b5",
X"1e",
X"c9",
X"06",
X"90",
X"2e",
X"b5",
X"16",
X"c9",
X"05",
X"f0",
X"27",
X"b9",
X"1e",
X"00",
X"0a",
X"90",
X"0a",
X"a9",
X"06",
X"20",
X"11",
X"da",
X"20",
X"95",
X"d7",
X"a4",
X"01",
X"98",
X"aa",
X"20",
X"95",
X"d7",
X"a6",
X"08",
X"bd",
X"25",
X"01",
X"18",
X"69",
X"04",
X"a6",
X"01",
X"20",
X"11",
X"da",
X"a6",
X"08",
X"fe",
X"25",
X"01",
X"60",
X"b9",
X"1e",
X"00",
X"c9",
X"06",
X"90",
X"1d",
X"b9",
X"16",
X"00",
X"c9",
X"05",
X"f0",
X"f1",
X"20",
X"95",
X"d7",
X"a4",
X"01",
X"b9",
X"25",
X"01",
X"18",
X"69",
X"04",
X"a6",
X"08",
X"20",
X"11",
X"da",
X"a6",
X"01",
X"fe",
X"25",
X"01",
X"60",
X"98",
X"aa",
X"20",
X"1c",
X"db",
X"a6",
X"08",
X"b5",
X"16",
X"c9",
X"0d",
X"f0",
X"22",
X"c9",
X"11",
X"f0",
X"1e",
X"c9",
X"05",
X"f0",
X"1a",
X"c9",
X"12",
X"f0",
X"08",
X"c9",
X"0e",
X"f0",
X"04",
X"c9",
X"07",
X"b0",
X"0e",
X"b5",
X"58",
X"49",
X"ff",
X"a8",
X"c8",
X"94",
X"58",
X"b5",
X"46",
X"49",
X"03",
X"95",
X"46",
X"60",
X"a9",
X"ff",
X"9d",
X"a2",
X"03",
X"ad",
X"47",
X"07",
X"d0",
X"29",
X"b5",
X"1e",
X"30",
X"25",
X"b5",
X"16",
X"c9",
X"24",
X"d0",
X"06",
X"b5",
X"1e",
X"aa",
X"20",
X"5f",
X"db",
X"20",
X"41",
X"dc",
X"b0",
X"14",
X"8a",
X"20",
X"54",
X"dc",
X"b5",
X"cf",
X"85",
X"00",
X"8a",
X"48",
X"20",
X"25",
X"e3",
X"68",
X"aa",
X"90",
X"03",
X"20",
X"bc",
X"db",
X"a6",
X"08",
X"60",
X"ad",
X"47",
X"07",
X"d0",
X"37",
X"9d",
X"a2",
X"03",
X"20",
X"41",
X"dc",
X"b0",
X"2f",
X"a9",
X"02",
X"85",
X"00",
X"a6",
X"08",
X"20",
X"52",
X"dc",
X"29",
X"02",
X"d0",
X"22",
X"b9",
X"ad",
X"04",
X"c9",
X"20",
X"90",
X"05",
X"20",
X"25",
X"e3",
X"b0",
X"19",
X"b9",
X"ad",
X"04",
X"18",
X"69",
X"80",
X"99",
X"ad",
X"04",
X"b9",
X"af",
X"04",
X"18",
X"69",
X"80",
X"99",
X"af",
X"04",
X"c6",
X"00",
X"d0",
X"d5",
X"a6",
X"08",
X"60",
X"a6",
X"08",
X"b9",
X"af",
X"04",
X"38",
X"ed",
X"ad",
X"04",
X"c9",
X"04",
X"b0",
X"08",
X"a5",
X"9f",
X"10",
X"04",
X"a9",
X"01",
X"85",
X"9f",
X"ad",
X"af",
X"04",
X"38",
X"f9",
X"ad",
X"04",
X"c9",
X"06",
X"b0",
X"1b",
X"a5",
X"9f",
X"30",
X"17",
X"a5",
X"00",
X"b4",
X"16",
X"c0",
X"2b",
X"f0",
X"05",
X"c0",
X"2c",
X"f0",
X"01",
X"8a",
X"a6",
X"08",
X"9d",
X"a2",
X"03",
X"a9",
X"00",
X"85",
X"1d",
X"60",
X"a9",
X"01",
X"85",
X"00",
X"ad",
X"ae",
X"04",
X"38",
X"f9",
X"ac",
X"04",
X"c9",
X"08",
X"90",
X"0d",
X"e6",
X"00",
X"b9",
X"ae",
X"04",
X"18",
X"ed",
X"ac",
X"04",
X"c9",
X"09",
X"b0",
X"03",
X"20",
X"4b",
X"df",
X"a6",
X"08",
X"60",
X"80",
X"00",
X"a8",
X"b5",
X"cf",
X"18",
X"79",
X"16",
X"dc",
X"2c",
X"b5",
X"cf",
X"a4",
X"0e",
X"c0",
X"0b",
X"f0",
X"17",
X"b4",
X"b6",
X"c0",
X"01",
X"d0",
X"11",
X"38",
X"e9",
X"20",
X"85",
X"ce",
X"98",
X"e9",
X"00",
X"85",
X"b5",
X"a9",
X"00",
X"85",
X"9f",
X"8d",
X"33",
X"04",
X"60",
X"ad",
X"d0",
X"03",
X"c9",
X"f0",
X"b0",
X"09",
X"a4",
X"b5",
X"88",
X"d0",
X"04",
X"a5",
X"ce",
X"c9",
X"d0",
X"60",
X"a5",
X"08",
X"0a",
X"0a",
X"18",
X"69",
X"04",
X"a8",
X"ad",
X"d1",
X"03",
X"29",
X"0f",
X"c9",
X"0f",
X"60",
X"20",
X"10",
X"ad",
X"16",
X"07",
X"d0",
X"2e",
X"a5",
X"0e",
X"c9",
X"0b",
X"f0",
X"28",
X"c9",
X"04",
X"90",
X"24",
X"a9",
X"01",
X"ac",
X"04",
X"07",
X"d0",
X"0a",
X"a5",
X"1d",
X"f0",
X"04",
X"c9",
X"03",
X"d0",
X"04",
X"a9",
X"02",
X"85",
X"1d",
X"a5",
X"b5",
X"c9",
X"01",
X"d0",
X"0b",
X"a9",
X"ff",
X"8d",
X"90",
X"04",
X"a5",
X"ce",
X"c9",
X"cf",
X"90",
X"01",
X"60",
X"a0",
X"02",
X"ad",
X"14",
X"07",
X"d0",
X"0c",
X"ad",
X"54",
X"07",
X"d0",
X"07",
X"88",
X"ad",
X"04",
X"07",
X"d0",
X"01",
X"88",
X"b9",
X"ad",
X"e3",
X"85",
X"eb",
X"a8",
X"ae",
X"54",
X"07",
X"ad",
X"14",
X"07",
X"f0",
X"01",
X"e8",
X"a5",
X"ce",
X"dd",
X"62",
X"dc",
X"90",
X"35",
X"20",
X"e9",
X"e3",
X"f0",
X"30",
X"20",
X"a1",
X"df",
X"b0",
X"4f",
X"a4",
X"9f",
X"10",
X"27",
X"a4",
X"04",
X"c0",
X"04",
X"90",
X"21",
X"20",
X"8f",
X"df",
X"b0",
X"10",
X"ac",
X"4e",
X"07",
X"f0",
X"13",
X"ac",
X"84",
X"07",
X"d0",
X"0e",
X"20",
X"ed",
X"bc",
X"4c",
X"f6",
X"dc",
X"c9",
X"26",
X"f0",
X"04",
X"a9",
X"02",
X"85",
X"ff",
X"a9",
X"01",
X"85",
X"9f",
X"a4",
X"eb",
X"a5",
X"ce",
X"c9",
X"cf",
X"b0",
X"60",
X"20",
X"e8",
X"e3",
X"20",
X"a1",
X"df",
X"b0",
X"14",
X"48",
X"20",
X"e8",
X"e3",
X"85",
X"00",
X"68",
X"85",
X"01",
X"d0",
X"0c",
X"a5",
X"00",
X"f0",
X"49",
X"20",
X"a1",
X"df",
X"90",
X"03",
X"4c",
X"05",
X"de",
X"20",
X"9a",
X"df",
X"b0",
X"3c",
X"a4",
X"9f",
X"30",
X"38",
X"c9",
X"c5",
X"d0",
X"03",
X"4c",
X"0e",
X"de",
X"20",
X"bd",
X"de",
X"f0",
X"2c",
X"ac",
X"0e",
X"07",
X"d0",
X"23",
X"a4",
X"04",
X"c0",
X"05",
X"90",
X"07",
X"a5",
X"45",
X"85",
X"00",
X"4c",
X"4b",
X"df",
X"20",
X"c4",
X"de",
X"a9",
X"f0",
X"25",
X"ce",
X"85",
X"ce",
X"20",
X"e8",
X"de",
X"a9",
X"00",
X"85",
X"9f",
X"8d",
X"33",
X"04",
X"8d",
X"84",
X"04",
X"a9",
X"00",
X"85",
X"1d",
X"a4",
X"eb",
X"c8",
X"c8",
X"a9",
X"02",
X"85",
X"00",
X"c8",
X"84",
X"eb",
X"a5",
X"ce",
X"c9",
X"20",
X"90",
X"16",
X"c9",
X"e4",
X"b0",
X"28",
X"20",
X"ec",
X"e3",
X"f0",
X"0d",
X"c9",
X"1c",
X"f0",
X"09",
X"c9",
X"6b",
X"f0",
X"05",
X"20",
X"9a",
X"df",
X"90",
X"17",
X"a4",
X"eb",
X"c8",
X"a5",
X"ce",
X"c9",
X"08",
X"90",
X"0d",
X"c9",
X"d0",
X"b0",
X"09",
X"20",
X"ec",
X"e3",
X"d0",
X"05",
X"c6",
X"00",
X"d0",
X"cb",
X"60",
X"20",
X"bd",
X"de",
X"f0",
X"61",
X"20",
X"9a",
X"df",
X"90",
X"03",
X"4c",
X"2e",
X"de",
X"20",
X"a1",
X"df",
X"b0",
X"57",
X"20",
X"dd",
X"de",
X"90",
X"08",
X"ad",
X"0e",
X"07",
X"d0",
X"4a",
X"4c",
X"ff",
X"dd",
X"a4",
X"1d",
X"c0",
X"00",
X"d0",
X"3e",
X"a4",
X"33",
X"88",
X"d0",
X"39",
X"c9",
X"6c",
X"f0",
X"04",
X"c9",
X"1f",
X"d0",
X"31",
X"ad",
X"c4",
X"03",
X"d0",
X"04",
X"a0",
X"10",
X"84",
X"ff",
X"09",
X"20",
X"8d",
X"c4",
X"03",
X"a5",
X"86",
X"29",
X"0f",
X"f0",
X"0e",
X"a0",
X"00",
X"ad",
X"1a",
X"07",
X"f0",
X"01",
X"c8",
X"b9",
X"03",
X"de",
X"8d",
X"de",
X"06",
X"a5",
X"0e",
X"c9",
X"07",
X"f0",
X"0c",
X"c9",
X"08",
X"d0",
X"08",
X"a9",
X"02",
X"85",
X"0e",
X"60",
X"20",
X"4b",
X"df",
X"60",
X"a0",
X"34",
X"20",
X"1c",
X"de",
X"ee",
X"48",
X"07",
X"4c",
X"fe",
X"bb",
X"a9",
X"00",
X"8d",
X"72",
X"07",
X"a9",
X"02",
X"8d",
X"70",
X"07",
X"a9",
X"18",
X"85",
X"57",
X"a4",
X"02",
X"a9",
X"00",
X"91",
X"06",
X"4c",
X"4d",
X"8a",
X"f9",
X"07",
X"ff",
X"00",
X"18",
X"22",
X"50",
X"68",
X"90",
X"a4",
X"04",
X"c0",
X"06",
X"90",
X"04",
X"c0",
X"0a",
X"90",
X"01",
X"60",
X"c9",
X"24",
X"f0",
X"04",
X"c9",
X"25",
X"d0",
X"39",
X"a5",
X"0e",
X"c9",
X"05",
X"f0",
X"41",
X"a9",
X"01",
X"85",
X"33",
X"ee",
X"23",
X"07",
X"a5",
X"0e",
X"c9",
X"04",
X"f0",
X"1f",
X"a9",
X"33",
X"20",
X"16",
X"97",
X"a9",
X"80",
X"85",
X"fc",
X"4a",
X"8d",
X"13",
X"07",
X"a2",
X"04",
X"a5",
X"ce",
X"8d",
X"0f",
X"07",
X"dd",
X"29",
X"de",
X"b0",
X"03",
X"ca",
X"d0",
X"f8",
X"8e",
X"0f",
X"01",
X"a9",
X"04",
X"85",
X"0e",
X"4c",
X"88",
X"de",
X"c9",
X"26",
X"d0",
X"0a",
X"a5",
X"ce",
X"c9",
X"20",
X"b0",
X"04",
X"a9",
X"01",
X"85",
X"0e",
X"a9",
X"03",
X"85",
X"1d",
X"a9",
X"00",
X"85",
X"57",
X"8d",
X"05",
X"07",
X"a5",
X"86",
X"38",
X"ed",
X"1c",
X"07",
X"c9",
X"10",
X"b0",
X"04",
X"a9",
X"02",
X"85",
X"33",
X"a4",
X"33",
X"a5",
X"06",
X"0a",
X"0a",
X"0a",
X"0a",
X"18",
X"79",
X"24",
X"de",
X"85",
X"86",
X"a5",
X"06",
X"d0",
X"09",
X"ad",
X"1b",
X"07",
X"18",
X"79",
X"26",
X"de",
X"85",
X"6d",
X"60",
X"c9",
X"5f",
X"f0",
X"02",
X"c9",
X"60",
X"60",
X"20",
X"dd",
X"de",
X"90",
X"13",
X"a9",
X"70",
X"8d",
X"09",
X"07",
X"a9",
X"f9",
X"8d",
X"db",
X"06",
X"a9",
X"03",
X"8d",
X"86",
X"07",
X"4a",
X"8d",
X"0e",
X"07",
X"60",
X"c9",
X"67",
X"f0",
X"05",
X"c9",
X"68",
X"18",
X"d0",
X"01",
X"38",
X"60",
X"a5",
X"0b",
X"29",
X"04",
X"f0",
X"5c",
X"a5",
X"00",
X"c9",
X"11",
X"d0",
X"56",
X"a5",
X"01",
X"c9",
X"10",
X"d0",
X"50",
X"a9",
X"30",
X"8d",
X"de",
X"06",
X"a9",
X"03",
X"85",
X"0e",
X"a9",
X"10",
X"85",
X"ff",
X"a9",
X"20",
X"8d",
X"c4",
X"03",
X"ad",
X"d6",
X"06",
X"f0",
X"39",
X"29",
X"03",
X"0a",
X"0a",
X"aa",
X"a5",
X"86",
X"c9",
X"60",
X"90",
X"06",
X"e8",
X"c9",
X"a0",
X"90",
X"01",
X"e8",
X"bc",
X"f2",
X"87",
X"88",
X"8c",
X"5f",
X"07",
X"be",
X"b4",
X"9c",
X"bd",
X"bc",
X"9c",
X"8d",
X"50",
X"07",
X"a9",
X"80",
X"85",
X"fc",
X"a9",
X"00",
X"8d",
X"51",
X"07",
X"8d",
X"60",
X"07",
X"8d",
X"5c",
X"07",
X"8d",
X"52",
X"07",
X"ee",
X"5d",
X"07",
X"ee",
X"57",
X"07",
X"60",
X"a9",
X"00",
X"a4",
X"57",
X"a6",
X"00",
X"ca",
X"d0",
X"0a",
X"e8",
X"c0",
X"00",
X"30",
X"28",
X"a9",
X"ff",
X"4c",
X"66",
X"df",
X"a2",
X"02",
X"c0",
X"01",
X"10",
X"1d",
X"a9",
X"01",
X"a0",
X"10",
X"8c",
X"85",
X"07",
X"a0",
X"00",
X"84",
X"57",
X"c9",
X"00",
X"10",
X"01",
X"88",
X"84",
X"00",
X"18",
X"65",
X"86",
X"85",
X"86",
X"a5",
X"6d",
X"65",
X"00",
X"85",
X"6d",
X"8a",
X"49",
X"ff",
X"2d",
X"90",
X"04",
X"8d",
X"90",
X"04",
X"60",
X"10",
X"61",
X"88",
X"c4",
X"20",
X"b0",
X"df",
X"dd",
X"8b",
X"df",
X"60",
X"24",
X"6d",
X"8a",
X"c6",
X"20",
X"b0",
X"df",
X"dd",
X"96",
X"df",
X"60",
X"c9",
X"c2",
X"f0",
X"06",
X"c9",
X"c3",
X"f0",
X"02",
X"18",
X"60",
X"a9",
X"01",
X"85",
X"fe",
X"60",
X"a8",
X"29",
X"c0",
X"0a",
X"2a",
X"2a",
X"aa",
X"98",
X"60",
X"01",
X"01",
X"02",
X"02",
X"02",
X"05",
X"10",
X"f0",
X"b5",
X"1e",
X"29",
X"20",
X"d0",
X"f1",
X"20",
X"5b",
X"e1",
X"90",
X"ec",
X"b4",
X"16",
X"c0",
X"12",
X"d0",
X"06",
X"b5",
X"cf",
X"c9",
X"25",
X"90",
X"e0",
X"c0",
X"0e",
X"d0",
X"03",
X"4c",
X"63",
X"e1",
X"c0",
X"05",
X"d0",
X"03",
X"4c",
X"85",
X"e1",
X"c0",
X"12",
X"f0",
X"08",
X"c0",
X"2e",
X"f0",
X"04",
X"c0",
X"07",
X"b0",
X"74",
X"20",
X"ae",
X"e1",
X"d0",
X"03",
X"4c",
X"e2",
X"e0",
X"20",
X"b5",
X"e1",
X"f0",
X"f8",
X"c9",
X"23",
X"d0",
X"64",
X"a4",
X"02",
X"a9",
X"00",
X"91",
X"06",
X"b5",
X"16",
X"c9",
X"15",
X"b0",
X"0c",
X"c9",
X"06",
X"d0",
X"03",
X"20",
X"8e",
X"e1",
X"a9",
X"01",
X"20",
X"11",
X"da",
X"c9",
X"09",
X"90",
X"10",
X"c9",
X"11",
X"b0",
X"0c",
X"c9",
X"0a",
X"90",
X"04",
X"c9",
X"0d",
X"90",
X"04",
X"29",
X"01",
X"95",
X"16",
X"b5",
X"1e",
X"29",
X"f0",
X"09",
X"02",
X"95",
X"1e",
X"d6",
X"cf",
X"d6",
X"cf",
X"b5",
X"16",
X"c9",
X"07",
X"f0",
X"07",
X"a9",
X"fd",
X"ac",
X"4e",
X"07",
X"d0",
X"02",
X"a9",
X"ff",
X"95",
X"a0",
X"a0",
X"01",
X"20",
X"43",
X"e1",
X"10",
X"01",
X"c8",
X"b5",
X"16",
X"c9",
X"33",
X"f0",
X"06",
X"c9",
X"08",
X"f0",
X"02",
X"94",
X"46",
X"88",
X"b9",
X"bf",
X"df",
X"95",
X"58",
X"60",
X"a5",
X"04",
X"38",
X"e9",
X"08",
X"c9",
X"05",
X"b0",
X"72",
X"b5",
X"1e",
X"29",
X"40",
X"d0",
X"57",
X"b5",
X"1e",
X"0a",
X"90",
X"03",
X"4c",
X"fe",
X"e0",
X"b5",
X"1e",
X"f0",
X"f9",
X"c9",
X"05",
X"f0",
X"1f",
X"c9",
X"03",
X"b0",
X"1a",
X"b5",
X"1e",
X"c9",
X"02",
X"d0",
X"15",
X"a9",
X"10",
X"b4",
X"16",
X"c0",
X"12",
X"d0",
X"02",
X"a9",
X"00",
X"9d",
X"96",
X"07",
X"a9",
X"03",
X"95",
X"1e",
X"20",
X"4f",
X"e1",
X"60",
X"b5",
X"16",
X"c9",
X"06",
X"f0",
X"22",
X"c9",
X"12",
X"d0",
X"0e",
X"a9",
X"01",
X"95",
X"46",
X"a9",
X"08",
X"95",
X"58",
X"a5",
X"09",
X"29",
X"07",
X"f0",
X"10",
X"a0",
X"01",
X"20",
X"43",
X"e1",
X"10",
X"01",
X"c8",
X"98",
X"d5",
X"46",
X"d0",
X"03",
X"20",
X"24",
X"e1",
X"20",
X"4f",
X"e1",
X"b5",
X"1e",
X"29",
X"80",
X"d0",
X"05",
X"a9",
X"00",
X"95",
X"1e",
X"60",
X"b5",
X"1e",
X"29",
X"bf",
X"95",
X"1e",
X"60",
X"b5",
X"16",
X"c9",
X"03",
X"d0",
X"04",
X"b5",
X"1e",
X"f0",
X"38",
X"b5",
X"1e",
X"a8",
X"0a",
X"90",
X"07",
X"b5",
X"1e",
X"09",
X"40",
X"4c",
X"fc",
X"e0",
X"b9",
X"b9",
X"df",
X"95",
X"1e",
X"b5",
X"cf",
X"c9",
X"20",
X"90",
X"1f",
X"a0",
X"16",
X"a9",
X"02",
X"85",
X"eb",
X"a5",
X"eb",
X"d5",
X"46",
X"d0",
X"0c",
X"a9",
X"01",
X"20",
X"88",
X"e3",
X"f0",
X"05",
X"20",
X"b5",
X"e1",
X"d0",
X"08",
X"c6",
X"eb",
X"c8",
X"c0",
X"18",
X"90",
X"e7",
X"60",
X"e0",
X"05",
X"f0",
X"09",
X"b5",
X"1e",
X"0a",
X"90",
X"04",
X"a9",
X"02",
X"85",
X"ff",
X"b5",
X"16",
X"c9",
X"05",
X"d0",
X"09",
X"a9",
X"00",
X"85",
X"00",
X"a0",
X"fa",
X"4c",
X"37",
X"ca",
X"4c",
X"36",
X"db",
X"b5",
X"87",
X"38",
X"e5",
X"86",
X"85",
X"00",
X"b5",
X"6e",
X"e5",
X"6d",
X"60",
X"20",
X"63",
X"c3",
X"b5",
X"cf",
X"29",
X"f0",
X"09",
X"08",
X"95",
X"cf",
X"60",
X"b5",
X"cf",
X"18",
X"69",
X"3e",
X"c9",
X"44",
X"60",
X"20",
X"5b",
X"e1",
X"90",
X"1a",
X"b5",
X"a0",
X"18",
X"69",
X"02",
X"c9",
X"03",
X"90",
X"11",
X"20",
X"ae",
X"e1",
X"f0",
X"0c",
X"20",
X"b5",
X"e1",
X"f0",
X"07",
X"20",
X"4f",
X"e1",
X"a9",
X"fd",
X"95",
X"a0",
X"4c",
X"fe",
X"e0",
X"20",
X"ae",
X"e1",
X"f0",
X"1d",
X"c9",
X"23",
X"d0",
X"08",
X"20",
X"95",
X"d7",
X"a9",
X"fc",
X"95",
X"a0",
X"60",
X"bd",
X"8a",
X"07",
X"d0",
X"0c",
X"b5",
X"1e",
X"29",
X"88",
X"95",
X"1e",
X"20",
X"4f",
X"e1",
X"4c",
X"fe",
X"e0",
X"b5",
X"1e",
X"09",
X"01",
X"95",
X"1e",
X"60",
X"a9",
X"00",
X"a0",
X"15",
X"4c",
X"88",
X"e3",
X"c9",
X"26",
X"f0",
X"0e",
X"c9",
X"c2",
X"f0",
X"0a",
X"c9",
X"c3",
X"f0",
X"06",
X"c9",
X"5f",
X"f0",
X"02",
X"c9",
X"60",
X"60",
X"b5",
X"d5",
X"c9",
X"18",
X"90",
X"21",
X"20",
X"9c",
X"e3",
X"f0",
X"1c",
X"20",
X"b5",
X"e1",
X"f0",
X"17",
X"b5",
X"a6",
X"30",
X"18",
X"b5",
X"3a",
X"d0",
X"14",
X"a9",
X"fd",
X"95",
X"a6",
X"a9",
X"01",
X"95",
X"3a",
X"b5",
X"d5",
X"29",
X"f8",
X"95",
X"d5",
X"60",
X"a9",
X"00",
X"95",
X"3a",
X"60",
X"a9",
X"80",
X"95",
X"24",
X"a9",
X"02",
X"85",
X"ff",
X"60",
X"02",
X"08",
X"0e",
X"20",
X"03",
X"14",
X"0d",
X"20",
X"02",
X"14",
X"0e",
X"20",
X"02",
X"09",
X"0e",
X"15",
X"00",
X"00",
X"18",
X"06",
X"00",
X"00",
X"20",
X"0d",
X"00",
X"00",
X"30",
X"0d",
X"00",
X"00",
X"08",
X"08",
X"06",
X"04",
X"0a",
X"08",
X"03",
X"0e",
X"0d",
X"14",
X"00",
X"02",
X"10",
X"15",
X"04",
X"04",
X"0c",
X"1c",
X"8a",
X"18",
X"69",
X"07",
X"aa",
X"a0",
X"02",
X"d0",
X"07",
X"8a",
X"18",
X"69",
X"09",
X"aa",
X"a0",
X"06",
X"20",
X"9c",
X"e2",
X"4c",
X"de",
X"e2",
X"a0",
X"48",
X"84",
X"00",
X"a0",
X"44",
X"4c",
X"52",
X"e2",
X"a0",
X"08",
X"84",
X"00",
X"a0",
X"04",
X"b5",
X"87",
X"38",
X"ed",
X"1c",
X"07",
X"85",
X"01",
X"b5",
X"6e",
X"ed",
X"1a",
X"07",
X"30",
X"06",
X"05",
X"01",
X"f0",
X"02",
X"a4",
X"00",
X"98",
X"2d",
X"d1",
X"03",
X"9d",
X"d8",
X"03",
X"d0",
X"19",
X"4c",
X"7c",
X"e2",
X"e8",
X"20",
X"f6",
X"f1",
X"ca",
X"c9",
X"fe",
X"b0",
X"0d",
X"8a",
X"18",
X"69",
X"01",
X"aa",
X"a0",
X"01",
X"20",
X"9c",
X"e2",
X"4c",
X"de",
X"e2",
X"8a",
X"0a",
X"0a",
X"a8",
X"a9",
X"ff",
X"99",
X"b0",
X"04",
X"99",
X"b1",
X"04",
X"99",
X"b2",
X"04",
X"99",
X"b3",
X"04",
X"60",
X"86",
X"00",
X"b9",
X"b8",
X"03",
X"85",
X"02",
X"b9",
X"ad",
X"03",
X"85",
X"01",
X"8a",
X"0a",
X"0a",
X"48",
X"a8",
X"bd",
X"99",
X"04",
X"0a",
X"0a",
X"aa",
X"a5",
X"01",
X"18",
X"7d",
X"fd",
X"e1",
X"99",
X"ac",
X"04",
X"a5",
X"01",
X"18",
X"7d",
X"ff",
X"e1",
X"99",
X"ae",
X"04",
X"e8",
X"c8",
X"a5",
X"02",
X"18",
X"7d",
X"fd",
X"e1",
X"99",
X"ac",
X"04",
X"a5",
X"02",
X"18",
X"7d",
X"ff",
X"e1",
X"99",
X"ae",
X"04",
X"68",
X"a8",
X"a6",
X"00",
X"60",
X"ad",
X"1c",
X"07",
X"18",
X"69",
X"80",
X"85",
X"02",
X"ad",
X"1a",
X"07",
X"69",
X"00",
X"85",
X"01",
X"b5",
X"86",
X"c5",
X"02",
X"b5",
X"6d",
X"e5",
X"01",
X"90",
X"15",
X"b9",
X"ae",
X"04",
X"30",
X"0d",
X"a9",
X"ff",
X"be",
X"ac",
X"04",
X"30",
X"03",
X"99",
X"ac",
X"04",
X"99",
X"ae",
X"04",
X"a6",
X"08",
X"60",
X"b9",
X"ac",
X"04",
X"10",
X"11",
X"c9",
X"a0",
X"90",
X"0d",
X"a9",
X"00",
X"be",
X"ae",
X"04",
X"10",
X"03",
X"99",
X"ae",
X"04",
X"99",
X"ac",
X"04",
X"a6",
X"08",
X"60",
X"a2",
X"00",
X"84",
X"06",
X"a9",
X"01",
X"85",
X"07",
X"b9",
X"ac",
X"04",
X"dd",
X"ac",
X"04",
X"b0",
X"2a",
X"dd",
X"ae",
X"04",
X"90",
X"12",
X"f0",
X"42",
X"b9",
X"ae",
X"04",
X"d9",
X"ac",
X"04",
X"90",
X"3a",
X"dd",
X"ac",
X"04",
X"b0",
X"35",
X"a4",
X"06",
X"60",
X"bd",
X"ae",
X"04",
X"dd",
X"ac",
X"04",
X"90",
X"2a",
X"b9",
X"ae",
X"04",
X"dd",
X"ac",
X"04",
X"b0",
X"22",
X"a4",
X"06",
X"60",
X"dd",
X"ac",
X"04",
X"f0",
X"1a",
X"dd",
X"ae",
X"04",
X"90",
X"15",
X"f0",
X"13",
X"d9",
X"ae",
X"04",
X"90",
X"0a",
X"f0",
X"08",
X"b9",
X"ae",
X"04",
X"dd",
X"ac",
X"04",
X"b0",
X"04",
X"18",
X"a4",
X"06",
X"60",
X"e8",
X"c8",
X"c6",
X"07",
X"10",
X"a9",
X"38",
X"a4",
X"06",
X"60",
X"48",
X"8a",
X"18",
X"69",
X"01",
X"aa",
X"68",
X"4c",
X"a5",
X"e3",
X"8a",
X"18",
X"69",
X"0d",
X"aa",
X"a0",
X"1b",
X"4c",
X"a3",
X"e3",
X"a0",
X"1a",
X"8a",
X"18",
X"69",
X"07",
X"aa",
X"a9",
X"00",
X"20",
X"f0",
X"e3",
X"a6",
X"08",
X"c9",
X"00",
X"60",
X"00",
X"07",
X"0e",
X"08",
X"03",
X"0c",
X"02",
X"02",
X"0d",
X"0d",
X"08",
X"03",
X"0c",
X"02",
X"02",
X"0d",
X"0d",
X"08",
X"03",
X"0c",
X"02",
X"02",
X"0d",
X"0d",
X"08",
X"00",
X"10",
X"04",
X"14",
X"04",
X"04",
X"04",
X"20",
X"20",
X"08",
X"18",
X"08",
X"18",
X"02",
X"20",
X"20",
X"08",
X"18",
X"08",
X"18",
X"12",
X"20",
X"20",
X"18",
X"18",
X"18",
X"18",
X"18",
X"14",
X"14",
X"06",
X"06",
X"08",
X"10",
X"c8",
X"a9",
X"00",
X"2c",
X"a9",
X"01",
X"a2",
X"00",
X"48",
X"84",
X"04",
X"b9",
X"b0",
X"e3",
X"18",
X"75",
X"86",
X"85",
X"05",
X"b5",
X"6d",
X"69",
X"00",
X"29",
X"01",
X"4a",
X"05",
X"05",
X"6a",
X"4a",
X"4a",
X"4a",
X"20",
X"e1",
X"9b",
X"a4",
X"04",
X"b5",
X"ce",
X"18",
X"79",
X"cc",
X"e3",
X"29",
X"f0",
X"38",
X"e9",
X"20",
X"85",
X"02",
X"a8",
X"b1",
X"06",
X"85",
X"03",
X"a4",
X"04",
X"68",
X"d0",
X"05",
X"b5",
X"ce",
X"4c",
X"2b",
X"e4",
X"b5",
X"86",
X"29",
X"0f",
X"85",
X"04",
X"a5",
X"03",
X"60",
X"ff",
X"00",
X"30",
X"84",
X"00",
X"ad",
X"b9",
X"03",
X"18",
X"79",
X"33",
X"e4",
X"be",
X"9a",
X"03",
X"bc",
X"e5",
X"06",
X"84",
X"02",
X"20",
X"ae",
X"e4",
X"ad",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"99",
X"0b",
X"02",
X"99",
X"13",
X"02",
X"18",
X"69",
X"06",
X"99",
X"07",
X"02",
X"99",
X"0f",
X"02",
X"99",
X"17",
X"02",
X"a9",
X"21",
X"99",
X"02",
X"02",
X"99",
X"0a",
X"02",
X"99",
X"12",
X"02",
X"09",
X"40",
X"99",
X"06",
X"02",
X"99",
X"0e",
X"02",
X"99",
X"16",
X"02",
X"a2",
X"05",
X"a9",
X"e1",
X"99",
X"01",
X"02",
X"c8",
X"c8",
X"c8",
X"c8",
X"ca",
X"10",
X"f4",
X"a4",
X"02",
X"a5",
X"00",
X"d0",
X"05",
X"a9",
X"e0",
X"99",
X"01",
X"02",
X"a2",
X"00",
X"ad",
X"9d",
X"03",
X"38",
X"f9",
X"00",
X"02",
X"c9",
X"64",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"c8",
X"c8",
X"c8",
X"c8",
X"e8",
X"e0",
X"06",
X"d0",
X"e7",
X"a4",
X"00",
X"60",
X"a2",
X"06",
X"99",
X"00",
X"02",
X"18",
X"69",
X"08",
X"c8",
X"c8",
X"c8",
X"c8",
X"ca",
X"d0",
X"f3",
X"a4",
X"02",
X"60",
X"04",
X"00",
X"04",
X"00",
X"00",
X"04",
X"00",
X"04",
X"00",
X"08",
X"00",
X"08",
X"08",
X"00",
X"08",
X"00",
X"80",
X"82",
X"81",
X"83",
X"81",
X"83",
X"80",
X"82",
X"03",
X"03",
X"c3",
X"c3",
X"bc",
X"f3",
X"06",
X"ad",
X"47",
X"07",
X"d0",
X"08",
X"b5",
X"2a",
X"29",
X"7f",
X"c9",
X"01",
X"f0",
X"04",
X"a2",
X"00",
X"f0",
X"07",
X"a5",
X"09",
X"4a",
X"4a",
X"29",
X"03",
X"aa",
X"ad",
X"be",
X"03",
X"18",
X"7d",
X"c4",
X"e4",
X"99",
X"00",
X"02",
X"18",
X"7d",
X"cc",
X"e4",
X"99",
X"04",
X"02",
X"ad",
X"b3",
X"03",
X"18",
X"7d",
X"c0",
X"e4",
X"99",
X"03",
X"02",
X"18",
X"7d",
X"c8",
X"e4",
X"99",
X"07",
X"02",
X"bd",
X"d0",
X"e4",
X"99",
X"01",
X"02",
X"bd",
X"d4",
X"e4",
X"99",
X"05",
X"02",
X"bd",
X"d8",
X"e4",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"a6",
X"08",
X"ad",
X"d6",
X"03",
X"29",
X"fc",
X"f0",
X"09",
X"a9",
X"00",
X"95",
X"2a",
X"a9",
X"f8",
X"20",
X"c1",
X"e5",
X"60",
X"f9",
X"50",
X"f7",
X"50",
X"fa",
X"fb",
X"f8",
X"fb",
X"f6",
X"fb",
X"bc",
X"e5",
X"06",
X"ad",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"18",
X"69",
X"08",
X"99",
X"07",
X"02",
X"99",
X"0b",
X"02",
X"18",
X"69",
X"0c",
X"85",
X"05",
X"b5",
X"cf",
X"20",
X"c1",
X"e5",
X"69",
X"08",
X"99",
X"08",
X"02",
X"ad",
X"0d",
X"01",
X"85",
X"02",
X"a9",
X"01",
X"85",
X"03",
X"85",
X"04",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"99",
X"0a",
X"02",
X"a9",
X"7e",
X"99",
X"01",
X"02",
X"99",
X"09",
X"02",
X"a9",
X"7f",
X"99",
X"05",
X"02",
X"ad",
X"0f",
X"07",
X"f0",
X"15",
X"98",
X"18",
X"69",
X"0c",
X"a8",
X"ad",
X"0f",
X"01",
X"0a",
X"aa",
X"bd",
X"41",
X"e5",
X"85",
X"00",
X"bd",
X"42",
X"e5",
X"20",
X"b2",
X"eb",
X"a6",
X"08",
X"bc",
X"e5",
X"06",
X"ad",
X"d1",
X"03",
X"29",
X"0e",
X"f0",
X"14",
X"a9",
X"f8",
X"99",
X"14",
X"02",
X"99",
X"10",
X"02",
X"99",
X"0c",
X"02",
X"99",
X"08",
X"02",
X"99",
X"04",
X"02",
X"99",
X"00",
X"02",
X"60",
X"bc",
X"e5",
X"06",
X"84",
X"02",
X"c8",
X"c8",
X"c8",
X"ad",
X"ae",
X"03",
X"20",
X"ae",
X"e4",
X"a6",
X"08",
X"b5",
X"cf",
X"20",
X"bb",
X"e5",
X"ac",
X"4e",
X"07",
X"c0",
X"03",
X"f0",
X"05",
X"ac",
X"cc",
X"06",
X"f0",
X"02",
X"a9",
X"f8",
X"bc",
X"e5",
X"06",
X"99",
X"10",
X"02",
X"99",
X"14",
X"02",
X"a9",
X"5b",
X"ae",
X"43",
X"07",
X"f0",
X"02",
X"a9",
X"75",
X"a6",
X"08",
X"c8",
X"20",
X"b5",
X"e5",
X"a9",
X"02",
X"c8",
X"20",
X"b5",
X"e5",
X"e8",
X"20",
X"f6",
X"f1",
X"ca",
X"bc",
X"e5",
X"06",
X"0a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"68",
X"0a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"04",
X"02",
X"68",
X"0a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"08",
X"02",
X"68",
X"0a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"0c",
X"02",
X"68",
X"0a",
X"48",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"10",
X"02",
X"68",
X"0a",
X"90",
X"05",
X"a9",
X"f8",
X"99",
X"14",
X"02",
X"ad",
X"d1",
X"03",
X"0a",
X"90",
X"03",
X"20",
X"b3",
X"e5",
X"60",
X"a5",
X"09",
X"4a",
X"b0",
X"02",
X"d6",
X"db",
X"b5",
X"db",
X"20",
X"c1",
X"e5",
X"ad",
X"b3",
X"03",
X"99",
X"03",
X"02",
X"18",
X"69",
X"08",
X"99",
X"07",
X"02",
X"a9",
X"02",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"a9",
X"f7",
X"99",
X"01",
X"02",
X"a9",
X"fb",
X"99",
X"05",
X"02",
X"4c",
X"bd",
X"e6",
X"60",
X"61",
X"62",
X"63",
X"bc",
X"f3",
X"06",
X"b5",
X"2a",
X"c9",
X"02",
X"b0",
X"c6",
X"b5",
X"db",
X"99",
X"00",
X"02",
X"18",
X"69",
X"08",
X"99",
X"04",
X"02",
X"ad",
X"b3",
X"03",
X"99",
X"03",
X"02",
X"99",
X"07",
X"02",
X"a5",
X"09",
X"4a",
X"29",
X"03",
X"aa",
X"bd",
X"82",
X"e6",
X"c8",
X"20",
X"c1",
X"e5",
X"88",
X"a9",
X"02",
X"99",
X"02",
X"02",
X"a9",
X"82",
X"99",
X"06",
X"02",
X"a6",
X"08",
X"60",
X"76",
X"77",
X"78",
X"79",
X"d6",
X"d6",
X"d9",
X"d9",
X"8d",
X"8d",
X"e4",
X"e4",
X"76",
X"77",
X"78",
X"79",
X"02",
X"01",
X"02",
X"01",
X"ac",
X"ea",
X"06",
X"ad",
X"b9",
X"03",
X"18",
X"69",
X"08",
X"85",
X"02",
X"ad",
X"ae",
X"03",
X"85",
X"05",
X"a6",
X"39",
X"bd",
X"ce",
X"e6",
X"0d",
X"ca",
X"03",
X"85",
X"04",
X"8a",
X"48",
X"0a",
X"0a",
X"aa",
X"a9",
X"01",
X"85",
X"07",
X"85",
X"03",
X"bd",
X"be",
X"e6",
X"85",
X"00",
X"bd",
X"bf",
X"e6",
X"20",
X"b2",
X"eb",
X"c6",
X"07",
X"10",
X"f1",
X"ac",
X"ea",
X"06",
X"68",
X"f0",
X"2f",
X"c9",
X"03",
X"f0",
X"2b",
X"85",
X"00",
X"a5",
X"09",
X"4a",
X"29",
X"03",
X"0d",
X"ca",
X"03",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"a6",
X"00",
X"ca",
X"f0",
X"06",
X"99",
X"0a",
X"02",
X"99",
X"0e",
X"02",
X"b9",
X"06",
X"02",
X"09",
X"40",
X"99",
X"06",
X"02",
X"b9",
X"0e",
X"02",
X"09",
X"40",
X"99",
X"0e",
X"02",
X"4c",
X"64",
X"eb",
X"fc",
X"fc",
X"aa",
X"ab",
X"ac",
X"ad",
X"fc",
X"fc",
X"ae",
X"af",
X"b0",
X"b1",
X"fc",
X"a5",
X"a6",
X"a7",
X"a8",
X"a9",
X"fc",
X"a0",
X"a1",
X"a2",
X"a3",
X"a4",
X"69",
X"a5",
X"6a",
X"a7",
X"a8",
X"a9",
X"6b",
X"a0",
X"6c",
X"a2",
X"a3",
X"a4",
X"fc",
X"fc",
X"96",
X"97",
X"98",
X"99",
X"fc",
X"fc",
X"9a",
X"9b",
X"9c",
X"9d",
X"fc",
X"fc",
X"8f",
X"8e",
X"8e",
X"8f",
X"fc",
X"fc",
X"95",
X"94",
X"94",
X"95",
X"fc",
X"fc",
X"dc",
X"dc",
X"df",
X"df",
X"dc",
X"dc",
X"dd",
X"dd",
X"de",
X"de",
X"fc",
X"fc",
X"b2",
X"b3",
X"b4",
X"b5",
X"fc",
X"fc",
X"b6",
X"b3",
X"b7",
X"b5",
X"fc",
X"fc",
X"70",
X"71",
X"72",
X"73",
X"fc",
X"fc",
X"6e",
X"6e",
X"6f",
X"6f",
X"fc",
X"fc",
X"6d",
X"6d",
X"6f",
X"6f",
X"fc",
X"fc",
X"6f",
X"6f",
X"6e",
X"6e",
X"fc",
X"fc",
X"6f",
X"6f",
X"6d",
X"6d",
X"fc",
X"fc",
X"f4",
X"f4",
X"f5",
X"f5",
X"fc",
X"fc",
X"f4",
X"f4",
X"f5",
X"f5",
X"fc",
X"fc",
X"f5",
X"f5",
X"f4",
X"f4",
X"fc",
X"fc",
X"f5",
X"f5",
X"f4",
X"f4",
X"fc",
X"fc",
X"fc",
X"fc",
X"ef",
X"ef",
X"b9",
X"b8",
X"bb",
X"ba",
X"bc",
X"bc",
X"fc",
X"fc",
X"bd",
X"bd",
X"bc",
X"bc",
X"7a",
X"7b",
X"da",
X"db",
X"d8",
X"d8",
X"cd",
X"cd",
X"ce",
X"ce",
X"cf",
X"cf",
X"7d",
X"7c",
X"d1",
X"8c",
X"d3",
X"d2",
X"7d",
X"7c",
X"89",
X"88",
X"8b",
X"8a",
X"d5",
X"d4",
X"e3",
X"e2",
X"d3",
X"d2",
X"d5",
X"d4",
X"e3",
X"e2",
X"8b",
X"8a",
X"e5",
X"e5",
X"e6",
X"e6",
X"eb",
X"eb",
X"ec",
X"ec",
X"ed",
X"ed",
X"ee",
X"ee",
X"fc",
X"fc",
X"d0",
X"d0",
X"d7",
X"d7",
X"bf",
X"be",
X"c1",
X"c0",
X"c2",
X"fc",
X"c4",
X"c3",
X"c6",
X"c5",
X"c8",
X"c7",
X"bf",
X"be",
X"ca",
X"c9",
X"c2",
X"fc",
X"c4",
X"c3",
X"c6",
X"c5",
X"cc",
X"cb",
X"fc",
X"fc",
X"e8",
X"e7",
X"ea",
X"e9",
X"f2",
X"f2",
X"f3",
X"f3",
X"f2",
X"f2",
X"f1",
X"f1",
X"f1",
X"f1",
X"fc",
X"fc",
X"f0",
X"f0",
X"fc",
X"fc",
X"fc",
X"fc",
X"0c",
X"0c",
X"00",
X"0c",
X"0c",
X"a8",
X"54",
X"3c",
X"ea",
X"18",
X"48",
X"48",
X"cc",
X"c0",
X"18",
X"18",
X"18",
X"90",
X"24",
X"ff",
X"48",
X"9c",
X"d2",
X"d8",
X"f0",
X"f6",
X"fc",
X"01",
X"02",
X"03",
X"02",
X"01",
X"01",
X"03",
X"03",
X"03",
X"01",
X"01",
X"02",
X"02",
X"21",
X"01",
X"02",
X"01",
X"01",
X"02",
X"ff",
X"02",
X"02",
X"01",
X"01",
X"02",
X"02",
X"02",
X"08",
X"18",
X"18",
X"19",
X"1a",
X"19",
X"18",
X"b5",
X"cf",
X"85",
X"02",
X"ad",
X"ae",
X"03",
X"85",
X"05",
X"bc",
X"e5",
X"06",
X"84",
X"eb",
X"a9",
X"00",
X"8d",
X"09",
X"01",
X"b5",
X"46",
X"85",
X"03",
X"bd",
X"c5",
X"03",
X"85",
X"04",
X"b5",
X"16",
X"c9",
X"0d",
X"d0",
X"0a",
X"b4",
X"58",
X"30",
X"06",
X"bc",
X"8a",
X"07",
X"f0",
X"01",
X"60",
X"b5",
X"1e",
X"85",
X"ed",
X"29",
X"1f",
X"a8",
X"b5",
X"16",
X"c9",
X"35",
X"d0",
X"08",
X"a0",
X"00",
X"a9",
X"01",
X"85",
X"03",
X"a9",
X"15",
X"c9",
X"33",
X"d0",
X"13",
X"c6",
X"02",
X"a9",
X"03",
X"bc",
X"8a",
X"07",
X"f0",
X"02",
X"09",
X"20",
X"85",
X"04",
X"a0",
X"00",
X"84",
X"ed",
X"a9",
X"08",
X"c9",
X"32",
X"d0",
X"08",
X"a0",
X"03",
X"ae",
X"0e",
X"07",
X"bd",
X"78",
X"e8",
X"85",
X"ef",
X"84",
X"ec",
X"a6",
X"08",
X"c9",
X"0c",
X"d0",
X"07",
X"b5",
X"a0",
X"30",
X"03",
X"ee",
X"09",
X"01",
X"ad",
X"6a",
X"03",
X"f0",
X"09",
X"a0",
X"16",
X"c9",
X"01",
X"f0",
X"01",
X"c8",
X"84",
X"ef",
X"a4",
X"ef",
X"c0",
X"06",
X"d0",
X"1d",
X"b5",
X"1e",
X"c9",
X"02",
X"90",
X"04",
X"a2",
X"04",
X"86",
X"ec",
X"29",
X"20",
X"0d",
X"47",
X"07",
X"d0",
X"0c",
X"a5",
X"09",
X"29",
X"08",
X"d0",
X"06",
X"a5",
X"03",
X"49",
X"03",
X"85",
X"03",
X"b9",
X"5b",
X"e8",
X"05",
X"04",
X"85",
X"04",
X"b9",
X"40",
X"e8",
X"aa",
X"a4",
X"ec",
X"ad",
X"6a",
X"03",
X"f0",
X"30",
X"c9",
X"01",
X"d0",
X"13",
X"ad",
X"63",
X"03",
X"10",
X"02",
X"a2",
X"de",
X"a5",
X"ed",
X"29",
X"20",
X"f0",
X"03",
X"8e",
X"09",
X"01",
X"4c",
X"4b",
X"ea",
X"ad",
X"63",
X"03",
X"29",
X"01",
X"f0",
X"02",
X"a2",
X"e4",
X"a5",
X"ed",
X"29",
X"20",
X"f0",
X"ee",
X"a5",
X"02",
X"38",
X"e9",
X"10",
X"85",
X"02",
X"4c",
X"46",
X"e9",
X"e0",
X"24",
X"d0",
X"11",
X"c0",
X"05",
X"d0",
X"0a",
X"a2",
X"30",
X"a9",
X"02",
X"85",
X"03",
X"a9",
X"05",
X"85",
X"ec",
X"4c",
X"ca",
X"e9",
X"e0",
X"90",
X"d0",
X"12",
X"a5",
X"ed",
X"29",
X"20",
X"d0",
X"09",
X"ad",
X"8f",
X"07",
X"c9",
X"10",
X"b0",
X"02",
X"a2",
X"96",
X"4c",
X"37",
X"ea",
X"a5",
X"ef",
X"c9",
X"04",
X"b0",
X"10",
X"c0",
X"02",
X"90",
X"0c",
X"a2",
X"5a",
X"a4",
X"ef",
X"c0",
X"02",
X"d0",
X"04",
X"a2",
X"7e",
X"e6",
X"02",
X"a5",
X"ec",
X"c9",
X"04",
X"d0",
X"1e",
X"a2",
X"72",
X"e6",
X"02",
X"a4",
X"ef",
X"c0",
X"02",
X"f0",
X"04",
X"a2",
X"66",
X"e6",
X"02",
X"c0",
X"06",
X"d0",
X"0c",
X"a2",
X"54",
X"a5",
X"ed",
X"29",
X"20",
X"d0",
X"04",
X"a2",
X"8a",
X"c6",
X"02",
X"a4",
X"08",
X"a5",
X"ef",
X"c9",
X"05",
X"d0",
X"0c",
X"a5",
X"ed",
X"f0",
X"24",
X"29",
X"08",
X"f0",
X"5d",
X"a2",
X"b4",
X"d0",
X"1c",
X"e0",
X"48",
X"f0",
X"18",
X"b9",
X"96",
X"07",
X"c9",
X"05",
X"b0",
X"4e",
X"e0",
X"3c",
X"d0",
X"0d",
X"c9",
X"01",
X"f0",
X"46",
X"e6",
X"02",
X"e6",
X"02",
X"e6",
X"02",
X"4c",
X"29",
X"ea",
X"a5",
X"ef",
X"c9",
X"06",
X"f0",
X"37",
X"c9",
X"08",
X"f0",
X"33",
X"c9",
X"0c",
X"f0",
X"2f",
X"c9",
X"18",
X"b0",
X"2b",
X"a0",
X"00",
X"c9",
X"15",
X"d0",
X"10",
X"c8",
X"ad",
X"5f",
X"07",
X"c9",
X"07",
X"b0",
X"1d",
X"a2",
X"a2",
X"a9",
X"03",
X"85",
X"ec",
X"d0",
X"15",
X"a5",
X"09",
X"39",
X"76",
X"e8",
X"d0",
X"0e",
X"a5",
X"ed",
X"29",
X"a0",
X"0d",
X"47",
X"07",
X"d0",
X"05",
X"8a",
X"18",
X"69",
X"06",
X"aa",
X"a5",
X"ed",
X"29",
X"20",
X"f0",
X"0e",
X"a5",
X"ef",
X"c9",
X"04",
X"90",
X"08",
X"a0",
X"01",
X"8c",
X"09",
X"01",
X"88",
X"84",
X"ec",
X"a4",
X"eb",
X"20",
X"aa",
X"eb",
X"20",
X"aa",
X"eb",
X"20",
X"aa",
X"eb",
X"a6",
X"08",
X"bc",
X"e5",
X"06",
X"a5",
X"ef",
X"c9",
X"08",
X"d0",
X"03",
X"4c",
X"64",
X"eb",
X"ad",
X"09",
X"01",
X"f0",
X"3d",
X"b9",
X"02",
X"02",
X"09",
X"80",
X"c8",
X"c8",
X"20",
X"b5",
X"e5",
X"88",
X"88",
X"98",
X"aa",
X"a5",
X"ef",
X"c9",
X"05",
X"f0",
X"0d",
X"c9",
X"11",
X"f0",
X"09",
X"c9",
X"15",
X"b0",
X"05",
X"8a",
X"18",
X"69",
X"08",
X"aa",
X"bd",
X"01",
X"02",
X"48",
X"bd",
X"05",
X"02",
X"48",
X"b9",
X"11",
X"02",
X"9d",
X"01",
X"02",
X"b9",
X"15",
X"02",
X"9d",
X"05",
X"02",
X"68",
X"99",
X"15",
X"02",
X"68",
X"99",
X"11",
X"02",
X"ad",
X"6a",
X"03",
X"d0",
X"b6",
X"a5",
X"ef",
X"a6",
X"ec",
X"c9",
X"05",
X"d0",
X"03",
X"4c",
X"64",
X"eb",
X"c9",
X"07",
X"f0",
X"1d",
X"c9",
X"0d",
X"f0",
X"19",
X"c9",
X"0c",
X"f0",
X"15",
X"c9",
X"12",
X"d0",
X"04",
X"e0",
X"05",
X"d0",
X"48",
X"c9",
X"15",
X"d0",
X"05",
X"a9",
X"42",
X"99",
X"16",
X"02",
X"e0",
X"02",
X"90",
X"3b",
X"ad",
X"6a",
X"03",
X"d0",
X"36",
X"b9",
X"02",
X"02",
X"29",
X"a3",
X"99",
X"02",
X"02",
X"99",
X"0a",
X"02",
X"99",
X"12",
X"02",
X"09",
X"40",
X"e0",
X"05",
X"d0",
X"02",
X"09",
X"80",
X"99",
X"06",
X"02",
X"99",
X"0e",
X"02",
X"99",
X"16",
X"02",
X"e0",
X"04",
X"d0",
X"13",
X"b9",
X"0a",
X"02",
X"09",
X"80",
X"99",
X"0a",
X"02",
X"99",
X"12",
X"02",
X"09",
X"40",
X"99",
X"0e",
X"02",
X"99",
X"16",
X"02",
X"a5",
X"ef",
X"c9",
X"11",
X"d0",
X"36",
X"ad",
X"09",
X"01",
X"d0",
X"21",
X"b9",
X"12",
X"02",
X"29",
X"81",
X"99",
X"12",
X"02",
X"b9",
X"16",
X"02",
X"09",
X"41",
X"99",
X"16",
X"02",
X"ae",
X"8f",
X"07",
X"e0",
X"10",
X"b0",
X"30",
X"99",
X"0e",
X"02",
X"29",
X"81",
X"99",
X"0a",
X"02",
X"90",
X"26",
X"b9",
X"02",
X"02",
X"29",
X"81",
X"99",
X"02",
X"02",
X"b9",
X"06",
X"02",
X"09",
X"41",
X"99",
X"06",
X"02",
X"a5",
X"ef",
X"c9",
X"18",
X"90",
X"10",
X"a9",
X"82",
X"99",
X"0a",
X"02",
X"99",
X"12",
X"02",
X"09",
X"40",
X"99",
X"0e",
X"02",
X"99",
X"16",
X"02",
X"a6",
X"08",
X"ad",
X"d1",
X"03",
X"4a",
X"4a",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"04",
X"20",
X"c1",
X"eb",
X"68",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"00",
X"20",
X"c1",
X"eb",
X"68",
X"4a",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"10",
X"20",
X"b7",
X"eb",
X"68",
X"4a",
X"48",
X"90",
X"05",
X"a9",
X"08",
X"20",
X"b7",
X"eb",
X"68",
X"4a",
X"90",
X"12",
X"20",
X"b7",
X"eb",
X"b5",
X"16",
X"c9",
X"0c",
X"f0",
X"09",
X"b5",
X"b6",
X"c9",
X"02",
X"d0",
X"03",
X"20",
X"98",
X"c9",
X"60",
X"bd",
X"3e",
X"e7",
X"85",
X"00",
X"bd",
X"3f",
X"e7",
X"85",
X"01",
X"4c",
X"82",
X"f2",
X"18",
X"7d",
X"e5",
X"06",
X"a8",
X"a9",
X"f8",
X"4c",
X"c1",
X"e5",
X"18",
X"7d",
X"e5",
X"06",
X"a8",
X"20",
X"4a",
X"ec",
X"99",
X"10",
X"02",
X"60",
X"85",
X"85",
X"86",
X"86",
X"ad",
X"bc",
X"03",
X"85",
X"02",
X"ad",
X"b1",
X"03",
X"85",
X"05",
X"a9",
X"03",
X"85",
X"04",
X"4a",
X"85",
X"03",
X"bc",
X"ec",
X"06",
X"a2",
X"00",
X"bd",
X"cd",
X"eb",
X"85",
X"00",
X"bd",
X"ce",
X"eb",
X"20",
X"b2",
X"eb",
X"e0",
X"04",
X"d0",
X"f1",
X"a6",
X"08",
X"bc",
X"ec",
X"06",
X"ad",
X"4e",
X"07",
X"c9",
X"01",
X"f0",
X"08",
X"a9",
X"86",
X"99",
X"01",
X"02",
X"99",
X"05",
X"02",
X"bd",
X"e8",
X"03",
X"c9",
X"c4",
X"d0",
X"24",
X"a9",
X"87",
X"c8",
X"20",
X"bb",
X"e5",
X"88",
X"a9",
X"03",
X"ae",
X"4e",
X"07",
X"ca",
X"f0",
X"01",
X"4a",
X"a6",
X"08",
X"99",
X"02",
X"02",
X"09",
X"40",
X"99",
X"06",
X"02",
X"09",
X"80",
X"99",
X"0e",
X"02",
X"29",
X"83",
X"99",
X"0a",
X"02",
X"ad",
X"d4",
X"03",
X"48",
X"29",
X"04",
X"f0",
X"08",
X"a9",
X"f8",
X"99",
X"04",
X"02",
X"99",
X"0c",
X"02",
X"68",
X"29",
X"08",
X"f0",
X"08",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"99",
X"08",
X"02",
X"60",
X"a9",
X"02",
X"85",
X"00",
X"a9",
X"75",
X"a4",
X"0e",
X"c0",
X"05",
X"f0",
X"06",
X"a9",
X"03",
X"85",
X"00",
X"a9",
X"84",
X"bc",
X"ec",
X"06",
X"c8",
X"20",
X"bb",
X"e5",
X"a5",
X"09",
X"0a",
X"0a",
X"0a",
X"0a",
X"29",
X"c0",
X"05",
X"00",
X"c8",
X"20",
X"bb",
X"e5",
X"88",
X"88",
X"ad",
X"bc",
X"03",
X"20",
X"c1",
X"e5",
X"ad",
X"b1",
X"03",
X"99",
X"03",
X"02",
X"bd",
X"f1",
X"03",
X"38",
X"ed",
X"1c",
X"07",
X"85",
X"00",
X"38",
X"ed",
X"b1",
X"03",
X"65",
X"00",
X"69",
X"06",
X"99",
X"07",
X"02",
X"ad",
X"bd",
X"03",
X"99",
X"08",
X"02",
X"99",
X"0c",
X"02",
X"ad",
X"b2",
X"03",
X"99",
X"0b",
X"02",
X"a5",
X"00",
X"38",
X"ed",
X"b2",
X"03",
X"65",
X"00",
X"69",
X"06",
X"99",
X"0f",
X"02",
X"ad",
X"d4",
X"03",
X"20",
X"46",
X"ec",
X"ad",
X"d4",
X"03",
X"0a",
X"90",
X"05",
X"a9",
X"f8",
X"20",
X"c1",
X"e5",
X"a5",
X"00",
X"10",
X"10",
X"b9",
X"03",
X"02",
X"d9",
X"07",
X"02",
X"90",
X"08",
X"a9",
X"f8",
X"99",
X"04",
X"02",
X"99",
X"0c",
X"02",
X"60",
X"bc",
X"f1",
X"06",
X"ad",
X"ba",
X"03",
X"99",
X"00",
X"02",
X"ad",
X"af",
X"03",
X"99",
X"03",
X"02",
X"a5",
X"09",
X"4a",
X"4a",
X"48",
X"29",
X"01",
X"49",
X"64",
X"99",
X"01",
X"02",
X"68",
X"4a",
X"4a",
X"a9",
X"02",
X"90",
X"02",
X"09",
X"c0",
X"99",
X"02",
X"02",
X"60",
X"68",
X"67",
X"66",
X"bc",
X"ec",
X"06",
X"b5",
X"24",
X"f6",
X"24",
X"4a",
X"29",
X"07",
X"c9",
X"03",
X"b0",
X"4a",
X"aa",
X"bd",
X"06",
X"ed",
X"c8",
X"20",
X"bb",
X"e5",
X"88",
X"a6",
X"08",
X"ad",
X"ba",
X"03",
X"38",
X"e9",
X"04",
X"99",
X"00",
X"02",
X"99",
X"08",
X"02",
X"18",
X"69",
X"08",
X"99",
X"04",
X"02",
X"99",
X"0c",
X"02",
X"ad",
X"af",
X"03",
X"38",
X"e9",
X"04",
X"99",
X"03",
X"02",
X"99",
X"07",
X"02",
X"18",
X"69",
X"08",
X"99",
X"0b",
X"02",
X"99",
X"0f",
X"02",
X"a9",
X"02",
X"99",
X"02",
X"02",
X"a9",
X"82",
X"99",
X"06",
X"02",
X"a9",
X"42",
X"99",
X"0a",
X"02",
X"a9",
X"c2",
X"99",
X"0e",
X"02",
X"60",
X"a9",
X"00",
X"95",
X"24",
X"60",
X"bc",
X"e5",
X"06",
X"a9",
X"5b",
X"c8",
X"20",
X"b5",
X"e5",
X"c8",
X"a9",
X"02",
X"20",
X"b5",
X"e5",
X"88",
X"88",
X"ad",
X"ae",
X"03",
X"99",
X"03",
X"02",
X"99",
X"0f",
X"02",
X"18",
X"69",
X"08",
X"99",
X"07",
X"02",
X"99",
X"13",
X"02",
X"18",
X"69",
X"08",
X"99",
X"0b",
X"02",
X"99",
X"17",
X"02",
X"b5",
X"cf",
X"aa",
X"48",
X"e0",
X"20",
X"b0",
X"02",
X"a9",
X"f8",
X"20",
X"be",
X"e5",
X"68",
X"18",
X"69",
X"80",
X"aa",
X"e0",
X"20",
X"b0",
X"02",
X"a9",
X"f8",
X"99",
X"0c",
X"02",
X"99",
X"10",
X"02",
X"99",
X"14",
X"02",
X"ad",
X"d1",
X"03",
X"48",
X"29",
X"08",
X"f0",
X"08",
X"a9",
X"f8",
X"99",
X"00",
X"02",
X"99",
X"0c",
X"02",
X"68",
X"48",
X"29",
X"04",
X"f0",
X"08",
X"a9",
X"f8",
X"99",
X"04",
X"02",
X"99",
X"10",
X"02",
X"68",
X"29",
X"02",
X"f0",
X"08",
X"a9",
X"f8",
X"99",
X"08",
X"02",
X"99",
X"14",
X"02",
X"a6",
X"08",
X"60",
X"a4",
X"b5",
X"88",
X"d0",
X"20",
X"ad",
X"d3",
X"03",
X"29",
X"08",
X"d0",
X"19",
X"bc",
X"ee",
X"06",
X"ad",
X"b0",
X"03",
X"99",
X"03",
X"02",
X"ad",
X"bb",
X"03",
X"99",
X"00",
X"02",
X"a9",
X"74",
X"99",
X"01",
X"02",
X"a9",
X"02",
X"99",
X"02",
X"02",
X"60",
X"20",
X"28",
X"c8",
X"18",
X"00",
X"40",
X"50",
X"58",
X"80",
X"88",
X"b8",
X"78",
X"60",
X"a0",
X"b0",
X"b8",
X"00",
X"01",
X"02",
X"03",
X"04",
X"05",
X"06",
X"07",
X"08",
X"09",
X"0a",
X"0b",
X"0c",
X"0d",
X"0e",
X"0f",
X"10",
X"11",
X"12",
X"13",
X"14",
X"15",
X"16",
X"17",
X"18",
X"19",
X"1a",
X"1b",
X"1c",
X"1d",
X"1e",
X"1f",
X"20",
X"21",
X"22",
X"23",
X"24",
X"25",
X"26",
X"27",
X"08",
X"09",
X"28",
X"29",
X"2a",
X"2b",
X"2c",
X"2d",
X"08",
X"09",
X"0a",
X"0b",
X"0c",
X"30",
X"2c",
X"2d",
X"08",
X"09",
X"0a",
X"0b",
X"2e",
X"2f",
X"2c",
X"2d",
X"08",
X"09",
X"28",
X"29",
X"2a",
X"2b",
X"5c",
X"5d",
X"08",
X"09",
X"0a",
X"0b",
X"0c",
X"0d",
X"5e",
X"5f",
X"fc",
X"fc",
X"08",
X"09",
X"58",
X"59",
X"5a",
X"5a",
X"08",
X"09",
X"28",
X"29",
X"2a",
X"2b",
X"0e",
X"0f",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"33",
X"34",
X"35",
X"fc",
X"fc",
X"fc",
X"fc",
X"36",
X"37",
X"38",
X"39",
X"fc",
X"fc",
X"fc",
X"fc",
X"3a",
X"37",
X"3b",
X"3c",
X"fc",
X"fc",
X"fc",
X"fc",
X"3d",
X"3e",
X"3f",
X"40",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"41",
X"42",
X"43",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"33",
X"44",
X"45",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"33",
X"44",
X"47",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"33",
X"48",
X"49",
X"fc",
X"fc",
X"fc",
X"fc",
X"32",
X"33",
X"90",
X"91",
X"fc",
X"fc",
X"fc",
X"fc",
X"3a",
X"37",
X"92",
X"93",
X"fc",
X"fc",
X"fc",
X"fc",
X"9e",
X"9e",
X"9f",
X"9f",
X"fc",
X"fc",
X"fc",
X"fc",
X"3a",
X"37",
X"4f",
X"4f",
X"fc",
X"fc",
X"00",
X"01",
X"4c",
X"4d",
X"4e",
X"4e",
X"00",
X"01",
X"4c",
X"4d",
X"4a",
X"4a",
X"4b",
X"4b",
X"31",
X"46",
X"ad",
X"9e",
X"07",
X"f0",
X"05",
X"a5",
X"09",
X"4a",
X"b0",
X"40",
X"a5",
X"0e",
X"c9",
X"0b",
X"f0",
X"47",
X"ad",
X"0b",
X"07",
X"d0",
X"3c",
X"ac",
X"04",
X"07",
X"f0",
X"31",
X"a5",
X"1d",
X"c9",
X"00",
X"f0",
X"2b",
X"20",
X"34",
X"ef",
X"a5",
X"09",
X"29",
X"04",
X"d0",
X"21",
X"aa",
X"ac",
X"e4",
X"06",
X"a5",
X"33",
X"4a",
X"b0",
X"04",
X"c8",
X"c8",
X"c8",
X"c8",
X"ad",
X"54",
X"07",
X"f0",
X"09",
X"b9",
X"19",
X"02",
X"cd",
X"b5",
X"ee",
X"f0",
X"07",
X"e8",
X"bd",
X"e7",
X"ee",
X"99",
X"19",
X"02",
X"60",
X"20",
X"ec",
X"ef",
X"4c",
X"45",
X"ef",
X"20",
X"b0",
X"f0",
X"4c",
X"45",
X"ef",
X"a0",
X"0e",
X"b9",
X"07",
X"ee",
X"8d",
X"d5",
X"06",
X"a9",
X"04",
X"20",
X"be",
X"ef",
X"20",
X"e9",
X"f0",
X"ad",
X"11",
X"07",
X"f0",
X"25",
X"a0",
X"00",
X"ad",
X"81",
X"07",
X"cd",
X"11",
X"07",
X"8c",
X"11",
X"07",
X"b0",
X"18",
X"8d",
X"11",
X"07",
X"a0",
X"07",
X"b9",
X"07",
X"ee",
X"8d",
X"d5",
X"06",
X"a0",
X"04",
X"a5",
X"57",
X"05",
X"0c",
X"f0",
X"01",
X"88",
X"98",
X"20",
X"be",
X"ef",
X"ad",
X"d0",
X"03",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"00",
X"a2",
X"03",
X"ad",
X"e4",
X"06",
X"18",
X"69",
X"18",
X"a8",
X"a9",
X"f8",
X"46",
X"00",
X"90",
X"03",
X"20",
X"c1",
X"e5",
X"98",
X"38",
X"e9",
X"08",
X"a8",
X"ca",
X"10",
X"ef",
X"60",
X"58",
X"01",
X"00",
X"60",
X"ff",
X"04",
X"a2",
X"05",
X"bd",
X"9e",
X"ef",
X"95",
X"02",
X"ca",
X"10",
X"f8",
X"a2",
X"b8",
X"a0",
X"04",
X"20",
X"dc",
X"ef",
X"ad",
X"26",
X"02",
X"09",
X"40",
X"8d",
X"22",
X"02",
X"60",
X"85",
X"07",
X"ad",
X"ad",
X"03",
X"8d",
X"55",
X"07",
X"85",
X"05",
X"ad",
X"b8",
X"03",
X"85",
X"02",
X"a5",
X"33",
X"85",
X"03",
X"ad",
X"c4",
X"03",
X"85",
X"04",
X"ae",
X"d5",
X"06",
X"ac",
X"e4",
X"06",
X"bd",
X"17",
X"ee",
X"85",
X"00",
X"bd",
X"18",
X"ee",
X"20",
X"b2",
X"eb",
X"c6",
X"07",
X"d0",
X"f1",
X"60",
X"a5",
X"1d",
X"c9",
X"03",
X"f0",
X"52",
X"c9",
X"02",
X"f0",
X"3e",
X"c9",
X"01",
X"d0",
X"11",
X"ad",
X"04",
X"07",
X"d0",
X"51",
X"a0",
X"06",
X"ad",
X"14",
X"07",
X"d0",
X"22",
X"a0",
X"00",
X"4c",
X"28",
X"f0",
X"a0",
X"06",
X"ad",
X"14",
X"07",
X"d0",
X"16",
X"a0",
X"02",
X"a5",
X"57",
X"05",
X"0c",
X"f0",
X"0e",
X"ad",
X"00",
X"07",
X"c9",
X"09",
X"90",
X"1b",
X"a5",
X"45",
X"25",
X"33",
X"d0",
X"15",
X"c8",
X"20",
X"91",
X"f0",
X"a9",
X"00",
X"8d",
X"0d",
X"07",
X"b9",
X"07",
X"ee",
X"60",
X"a0",
X"04",
X"20",
X"91",
X"f0",
X"4c",
X"62",
X"f0",
X"a0",
X"04",
X"20",
X"91",
X"f0",
X"4c",
X"68",
X"f0",
X"a0",
X"05",
X"a5",
X"9f",
X"f0",
X"de",
X"20",
X"91",
X"f0",
X"4c",
X"6d",
X"f0",
X"a0",
X"01",
X"20",
X"91",
X"f0",
X"ad",
X"82",
X"07",
X"0d",
X"0d",
X"07",
X"d0",
X"0b",
X"a5",
X"0a",
X"0a",
X"b0",
X"06",
X"ad",
X"0d",
X"07",
X"4c",
X"d0",
X"f0",
X"a9",
X"03",
X"4c",
X"6f",
X"f0",
X"a9",
X"02",
X"85",
X"00",
X"20",
X"62",
X"f0",
X"48",
X"ad",
X"81",
X"07",
X"d0",
X"15",
X"ad",
X"0c",
X"07",
X"8d",
X"81",
X"07",
X"ad",
X"0d",
X"07",
X"18",
X"69",
X"01",
X"c5",
X"00",
X"90",
X"02",
X"a9",
X"00",
X"8d",
X"0d",
X"07",
X"68",
X"60",
X"ad",
X"54",
X"07",
X"f0",
X"05",
X"98",
X"18",
X"69",
X"08",
X"a8",
X"60",
X"00",
X"01",
X"00",
X"01",
X"00",
X"01",
X"02",
X"00",
X"01",
X"02",
X"02",
X"00",
X"02",
X"00",
X"02",
X"00",
X"02",
X"00",
X"02",
X"00",
X"ac",
X"0d",
X"07",
X"a5",
X"09",
X"29",
X"03",
X"d0",
X"0d",
X"c8",
X"c0",
X"0a",
X"90",
X"05",
X"a0",
X"00",
X"8c",
X"0b",
X"07",
X"8c",
X"0d",
X"07",
X"ad",
X"54",
X"07",
X"d0",
X"0c",
X"b9",
X"9c",
X"f0",
X"a0",
X"0f",
X"0a",
X"0a",
X"0a",
X"79",
X"07",
X"ee",
X"60",
X"98",
X"18",
X"69",
X"0a",
X"aa",
X"a0",
X"09",
X"bd",
X"9c",
X"f0",
X"d0",
X"02",
X"a0",
X"01",
X"b9",
X"07",
X"ee",
X"60",
X"ac",
X"e4",
X"06",
X"a5",
X"0e",
X"c9",
X"0b",
X"f0",
X"13",
X"ad",
X"d5",
X"06",
X"c9",
X"50",
X"f0",
X"1e",
X"c9",
X"b8",
X"f0",
X"1a",
X"c9",
X"c0",
X"f0",
X"16",
X"c9",
X"c8",
X"d0",
X"24",
X"b9",
X"12",
X"02",
X"29",
X"3f",
X"99",
X"12",
X"02",
X"b9",
X"16",
X"02",
X"29",
X"3f",
X"09",
X"40",
X"99",
X"16",
X"02",
X"b9",
X"1a",
X"02",
X"29",
X"3f",
X"99",
X"1a",
X"02",
X"b9",
X"1e",
X"02",
X"29",
X"3f",
X"09",
X"40",
X"99",
X"1e",
X"02",
X"60",
X"a2",
X"00",
X"a0",
X"00",
X"4c",
X"42",
X"f1",
X"a0",
X"01",
X"20",
X"a8",
X"f1",
X"a0",
X"03",
X"4c",
X"42",
X"f1",
X"a0",
X"00",
X"20",
X"a8",
X"f1",
X"a0",
X"02",
X"20",
X"71",
X"f1",
X"a6",
X"08",
X"60",
X"a0",
X"02",
X"20",
X"a8",
X"f1",
X"a0",
X"06",
X"4c",
X"42",
X"f1",
X"a9",
X"01",
X"a0",
X"01",
X"4c",
X"65",
X"f1",
X"a9",
X"09",
X"a0",
X"04",
X"20",
X"65",
X"f1",
X"e8",
X"e8",
X"a9",
X"09",
X"c8",
X"86",
X"00",
X"18",
X"65",
X"00",
X"aa",
X"20",
X"71",
X"f1",
X"a6",
X"08",
X"60",
X"b5",
X"ce",
X"99",
X"b8",
X"03",
X"b5",
X"86",
X"38",
X"ed",
X"1c",
X"07",
X"99",
X"ad",
X"03",
X"60",
X"a2",
X"00",
X"a0",
X"00",
X"4c",
X"c0",
X"f1",
X"a0",
X"00",
X"20",
X"a8",
X"f1",
X"a0",
X"02",
X"4c",
X"c0",
X"f1",
X"a0",
X"01",
X"20",
X"a8",
X"f1",
X"a0",
X"03",
X"4c",
X"c0",
X"f1",
X"a0",
X"02",
X"20",
X"a8",
X"f1",
X"a0",
X"06",
X"4c",
X"c0",
X"f1",
X"07",
X"16",
X"0d",
X"8a",
X"18",
X"79",
X"a5",
X"f1",
X"aa",
X"60",
X"a9",
X"01",
X"a0",
X"01",
X"4c",
X"ba",
X"f1",
X"a9",
X"09",
X"a0",
X"04",
X"86",
X"00",
X"18",
X"65",
X"00",
X"aa",
X"98",
X"48",
X"20",
X"d7",
X"f1",
X"0a",
X"0a",
X"0a",
X"0a",
X"05",
X"00",
X"85",
X"00",
X"68",
X"a8",
X"a5",
X"00",
X"99",
X"d0",
X"03",
X"a6",
X"08",
X"60",
X"20",
X"f6",
X"f1",
X"4a",
X"4a",
X"4a",
X"4a",
X"85",
X"00",
X"4c",
X"39",
X"f2",
X"7f",
X"3f",
X"1f",
X"0f",
X"07",
X"03",
X"01",
X"00",
X"80",
X"c0",
X"e0",
X"f0",
X"f8",
X"fc",
X"fe",
X"ff",
X"07",
X"0f",
X"07",
X"86",
X"04",
X"a0",
X"01",
X"b9",
X"1c",
X"07",
X"38",
X"f5",
X"86",
X"85",
X"07",
X"b9",
X"1a",
X"07",
X"f5",
X"6d",
X"be",
X"f3",
X"f1",
X"c9",
X"00",
X"30",
X"10",
X"be",
X"f4",
X"f1",
X"c9",
X"01",
X"10",
X"09",
X"a9",
X"38",
X"85",
X"06",
X"a9",
X"08",
X"20",
X"6d",
X"f2",
X"bd",
X"e3",
X"f1",
X"a6",
X"04",
X"c9",
X"00",
X"d0",
X"03",
X"88",
X"10",
X"d0",
X"60",
X"00",
X"08",
X"0c",
X"0e",
X"0f",
X"07",
X"03",
X"01",
X"00",
X"04",
X"00",
X"04",
X"ff",
X"00",
X"86",
X"04",
X"a0",
X"01",
X"b9",
X"37",
X"f2",
X"38",
X"f5",
X"ce",
X"85",
X"07",
X"a9",
X"01",
X"f5",
X"b5",
X"be",
X"34",
X"f2",
X"c9",
X"00",
X"30",
X"10",
X"be",
X"35",
X"f2",
X"c9",
X"01",
X"10",
X"09",
X"a9",
X"20",
X"85",
X"06",
X"a9",
X"04",
X"20",
X"6d",
X"f2",
X"bd",
X"2b",
X"f2",
X"a6",
X"04",
X"c9",
X"00",
X"d0",
X"03",
X"88",
X"10",
X"d1",
X"60",
X"85",
X"05",
X"a5",
X"07",
X"c5",
X"06",
X"b0",
X"0c",
X"4a",
X"4a",
X"4a",
X"29",
X"07",
X"c0",
X"01",
X"b0",
X"02",
X"65",
X"05",
X"aa",
X"60",
X"a5",
X"03",
X"4a",
X"4a",
X"a5",
X"00",
X"90",
X"0c",
X"99",
X"05",
X"02",
X"a5",
X"01",
X"99",
X"01",
X"02",
X"a9",
X"40",
X"d0",
X"0a",
X"99",
X"01",
X"02",
X"a5",
X"01",
X"99",
X"05",
X"02",
X"a9",
X"00",
X"05",
X"04",
X"99",
X"02",
X"02",
X"99",
X"06",
X"02",
X"a5",
X"02",
X"99",
X"00",
X"02",
X"99",
X"04",
X"02",
X"a5",
X"05",
X"99",
X"03",
X"02",
X"18",
X"69",
X"08",
X"99",
X"07",
X"02",
X"a5",
X"02",
X"18",
X"69",
X"08",
X"85",
X"02",
X"98",
X"18",
X"69",
X"08",
X"a8",
X"e8",
X"e8",
X"60",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ff",
X"ad",
X"70",
X"07",
X"d0",
X"04",
X"8d",
X"15",
X"40",
X"60",
X"a9",
X"ff",
X"8d",
X"17",
X"40",
X"a9",
X"0f",
X"8d",
X"15",
X"40",
X"ad",
X"c6",
X"07",
X"d0",
X"06",
X"a5",
X"fa",
X"c9",
X"01",
X"d0",
X"5d",
X"ad",
X"b2",
X"07",
X"d0",
X"23",
X"a5",
X"fa",
X"f0",
X"66",
X"8d",
X"b2",
X"07",
X"8d",
X"c6",
X"07",
X"a9",
X"00",
X"8d",
X"15",
X"40",
X"85",
X"f1",
X"85",
X"f2",
X"85",
X"f3",
X"a9",
X"0f",
X"8d",
X"15",
X"40",
X"a9",
X"2a",
X"8d",
X"bb",
X"07",
X"a9",
X"44",
X"d0",
X"11",
X"ad",
X"bb",
X"07",
X"c9",
X"24",
X"f0",
X"08",
X"c9",
X"1e",
X"f0",
X"f1",
X"c9",
X"18",
X"d0",
X"09",
X"a9",
X"64",
X"a2",
X"84",
X"a0",
X"7f",
X"20",
X"88",
X"f3",
X"ce",
X"bb",
X"07",
X"d0",
X"2a",
X"a9",
X"00",
X"8d",
X"15",
X"40",
X"ad",
X"b2",
X"07",
X"c9",
X"02",
X"d0",
X"05",
X"a9",
X"00",
X"8d",
X"c6",
X"07",
X"a9",
X"00",
X"8d",
X"b2",
X"07",
X"f0",
X"12",
X"20",
X"1b",
X"f4",
X"20",
X"7c",
X"f5",
X"20",
X"67",
X"f6",
X"20",
X"94",
X"f6",
X"a9",
X"00",
X"85",
X"fb",
X"85",
X"fc",
X"a9",
X"00",
X"85",
X"ff",
X"85",
X"fe",
X"85",
X"fd",
X"85",
X"fa",
X"ac",
X"c0",
X"07",
X"a5",
X"f4",
X"29",
X"03",
X"f0",
X"07",
X"ee",
X"c0",
X"07",
X"c0",
X"30",
X"90",
X"06",
X"98",
X"f0",
X"03",
X"ce",
X"c0",
X"07",
X"8c",
X"11",
X"40",
X"60",
X"8c",
X"01",
X"40",
X"8e",
X"00",
X"40",
X"60",
X"20",
X"81",
X"f3",
X"a2",
X"00",
X"a8",
X"b9",
X"01",
X"ff",
X"f0",
X"0b",
X"9d",
X"02",
X"40",
X"b9",
X"00",
X"ff",
X"09",
X"08",
X"9d",
X"03",
X"40",
X"60",
X"8e",
X"04",
X"40",
X"8c",
X"05",
X"40",
X"60",
X"20",
X"9f",
X"f3",
X"a2",
X"04",
X"d0",
X"e0",
X"a2",
X"08",
X"d0",
X"dc",
X"9f",
X"9b",
X"98",
X"96",
X"95",
X"94",
X"92",
X"90",
X"90",
X"9a",
X"97",
X"95",
X"93",
X"92",
X"a9",
X"40",
X"8d",
X"bb",
X"07",
X"a9",
X"62",
X"20",
X"8b",
X"f3",
X"a2",
X"99",
X"d0",
X"25",
X"a9",
X"26",
X"d0",
X"02",
X"a9",
X"18",
X"a2",
X"82",
X"a0",
X"a7",
X"20",
X"88",
X"f3",
X"a9",
X"28",
X"8d",
X"bb",
X"07",
X"ad",
X"bb",
X"07",
X"c9",
X"25",
X"d0",
X"06",
X"a2",
X"5f",
X"a0",
X"f6",
X"d0",
X"08",
X"c9",
X"20",
X"d0",
X"29",
X"a2",
X"48",
X"a0",
X"bc",
X"20",
X"81",
X"f3",
X"d0",
X"20",
X"a9",
X"05",
X"a0",
X"99",
X"d0",
X"04",
X"a9",
X"0a",
X"a0",
X"93",
X"a2",
X"9e",
X"8d",
X"bb",
X"07",
X"a9",
X"0c",
X"20",
X"88",
X"f3",
X"ad",
X"bb",
X"07",
X"c9",
X"06",
X"d0",
X"05",
X"a9",
X"bb",
X"8d",
X"01",
X"40",
X"d0",
X"60",
X"a4",
X"ff",
X"f0",
X"20",
X"84",
X"f1",
X"30",
X"aa",
X"46",
X"ff",
X"b0",
X"aa",
X"46",
X"ff",
X"b0",
X"d4",
X"46",
X"ff",
X"b0",
X"2c",
X"46",
X"ff",
X"b0",
X"4a",
X"46",
X"ff",
X"b0",
X"7f",
X"46",
X"ff",
X"b0",
X"be",
X"46",
X"ff",
X"b0",
X"80",
X"a5",
X"f1",
X"f0",
X"17",
X"30",
X"9a",
X"4a",
X"b0",
X"97",
X"4a",
X"b0",
X"c2",
X"4a",
X"b0",
X"1b",
X"4a",
X"b0",
X"3c",
X"4a",
X"b0",
X"67",
X"4a",
X"b0",
X"b6",
X"4a",
X"b0",
X"48",
X"60",
X"a9",
X"0e",
X"8d",
X"bb",
X"07",
X"a0",
X"9c",
X"a2",
X"9e",
X"a9",
X"26",
X"20",
X"88",
X"f3",
X"ac",
X"bb",
X"07",
X"b9",
X"b0",
X"f3",
X"8d",
X"00",
X"40",
X"c0",
X"06",
X"d0",
X"05",
X"a9",
X"9e",
X"8d",
X"02",
X"40",
X"d0",
X"25",
X"a9",
X"0e",
X"a0",
X"cb",
X"a2",
X"9f",
X"8d",
X"bb",
X"07",
X"a9",
X"28",
X"20",
X"88",
X"f3",
X"d0",
X"15",
X"ac",
X"bb",
X"07",
X"c0",
X"08",
X"d0",
X"09",
X"a9",
X"a0",
X"8d",
X"02",
X"40",
X"a9",
X"9f",
X"d0",
X"02",
X"a9",
X"90",
X"8d",
X"00",
X"40",
X"ce",
X"bb",
X"07",
X"d0",
X"0e",
X"a2",
X"00",
X"86",
X"f1",
X"a2",
X"0e",
X"8e",
X"15",
X"40",
X"a2",
X"0f",
X"8e",
X"15",
X"40",
X"60",
X"a9",
X"2f",
X"8d",
X"bb",
X"07",
X"ad",
X"bb",
X"07",
X"4a",
X"b0",
X"10",
X"4a",
X"b0",
X"0d",
X"29",
X"02",
X"f0",
X"09",
X"a0",
X"91",
X"a2",
X"9a",
X"a9",
X"44",
X"20",
X"88",
X"f3",
X"4c",
X"a2",
X"f4",
X"58",
X"02",
X"54",
X"56",
X"4e",
X"44",
X"4c",
X"52",
X"4c",
X"48",
X"3e",
X"36",
X"3e",
X"36",
X"30",
X"28",
X"4a",
X"50",
X"4a",
X"64",
X"3c",
X"32",
X"3c",
X"32",
X"2c",
X"24",
X"3a",
X"64",
X"3a",
X"34",
X"2c",
X"22",
X"2c",
X"22",
X"1c",
X"14",
X"14",
X"04",
X"22",
X"24",
X"16",
X"04",
X"24",
X"26",
X"18",
X"04",
X"26",
X"28",
X"1a",
X"04",
X"28",
X"2a",
X"1c",
X"04",
X"2a",
X"2c",
X"1e",
X"04",
X"2c",
X"2e",
X"20",
X"04",
X"2e",
X"30",
X"22",
X"04",
X"30",
X"32",
X"a9",
X"35",
X"a2",
X"8d",
X"d0",
X"04",
X"a9",
X"06",
X"a2",
X"98",
X"8d",
X"bd",
X"07",
X"a0",
X"7f",
X"a9",
X"42",
X"20",
X"a6",
X"f3",
X"ad",
X"bd",
X"07",
X"c9",
X"30",
X"d0",
X"05",
X"a9",
X"54",
X"8d",
X"06",
X"40",
X"d0",
X"2e",
X"a9",
X"20",
X"8d",
X"bd",
X"07",
X"a0",
X"94",
X"a9",
X"5e",
X"d0",
X"0b",
X"ad",
X"bd",
X"07",
X"c9",
X"18",
X"d0",
X"1c",
X"a0",
X"93",
X"a9",
X"18",
X"d0",
X"7f",
X"a9",
X"36",
X"8d",
X"bd",
X"07",
X"ad",
X"bd",
X"07",
X"4a",
X"b0",
X"0b",
X"a8",
X"b9",
X"d9",
X"f4",
X"a2",
X"5d",
X"a0",
X"7f",
X"20",
X"a6",
X"f3",
X"ce",
X"bd",
X"07",
X"d0",
X"0e",
X"a2",
X"00",
X"86",
X"f2",
X"a2",
X"0d",
X"8e",
X"15",
X"40",
X"a2",
X"0f",
X"8e",
X"15",
X"40",
X"60",
X"a5",
X"f2",
X"29",
X"40",
X"d0",
X"65",
X"a4",
X"fe",
X"f0",
X"20",
X"84",
X"f2",
X"30",
X"3e",
X"46",
X"fe",
X"b0",
X"8a",
X"46",
X"fe",
X"b0",
X"6a",
X"46",
X"fe",
X"b0",
X"6a",
X"46",
X"fe",
X"b0",
X"a0",
X"46",
X"fe",
X"b0",
X"80",
X"46",
X"fe",
X"b0",
X"b0",
X"46",
X"fe",
X"b0",
X"3c",
X"a5",
X"f2",
X"f0",
X"17",
X"30",
X"27",
X"4a",
X"b0",
X"13",
X"4a",
X"b0",
X"5d",
X"4a",
X"b0",
X"5a",
X"4a",
X"b0",
X"8d",
X"4a",
X"b0",
X"07",
X"4a",
X"b0",
X"99",
X"4a",
X"b0",
X"26",
X"60",
X"4c",
X"2c",
X"f5",
X"4c",
X"68",
X"f5",
X"a9",
X"38",
X"8d",
X"bd",
X"07",
X"a0",
X"c4",
X"a9",
X"18",
X"d0",
X"0b",
X"ad",
X"bd",
X"07",
X"c9",
X"08",
X"d0",
X"8e",
X"a0",
X"a4",
X"a9",
X"5a",
X"a2",
X"9f",
X"d0",
X"83",
X"a9",
X"30",
X"8d",
X"bd",
X"07",
X"ad",
X"bd",
X"07",
X"a2",
X"03",
X"4a",
X"b0",
X"d6",
X"ca",
X"d0",
X"fa",
X"a8",
X"b9",
X"d3",
X"f4",
X"a2",
X"82",
X"a0",
X"7f",
X"d0",
X"e4",
X"a9",
X"10",
X"d0",
X"02",
X"a9",
X"20",
X"8d",
X"bd",
X"07",
X"a9",
X"7f",
X"8d",
X"05",
X"40",
X"a9",
X"00",
X"8d",
X"be",
X"07",
X"ee",
X"be",
X"07",
X"ad",
X"be",
X"07",
X"4a",
X"a8",
X"cc",
X"bd",
X"07",
X"f0",
X"0c",
X"a9",
X"9d",
X"8d",
X"04",
X"40",
X"b9",
X"f8",
X"f4",
X"20",
X"a9",
X"f3",
X"60",
X"4c",
X"6d",
X"f5",
X"01",
X"0e",
X"0e",
X"0d",
X"0b",
X"06",
X"0c",
X"0f",
X"0a",
X"09",
X"03",
X"0d",
X"08",
X"0d",
X"06",
X"0c",
X"a9",
X"20",
X"8d",
X"bf",
X"07",
X"ad",
X"bf",
X"07",
X"4a",
X"90",
X"12",
X"a8",
X"be",
X"2b",
X"f6",
X"b9",
X"ea",
X"ff",
X"8d",
X"0c",
X"40",
X"8e",
X"0e",
X"40",
X"a9",
X"18",
X"8d",
X"0f",
X"40",
X"ce",
X"bf",
X"07",
X"d0",
X"09",
X"a9",
X"f0",
X"8d",
X"0c",
X"40",
X"a9",
X"00",
X"85",
X"f3",
X"60",
X"a4",
X"fd",
X"f0",
X"0a",
X"84",
X"f3",
X"46",
X"fd",
X"b0",
X"ca",
X"46",
X"fd",
X"b0",
X"0b",
X"a5",
X"f3",
X"f0",
X"06",
X"4a",
X"b0",
X"c4",
X"4a",
X"b0",
X"06",
X"60",
X"a9",
X"40",
X"8d",
X"bf",
X"07",
X"ad",
X"bf",
X"07",
X"4a",
X"a8",
X"a2",
X"0f",
X"b9",
X"c9",
X"ff",
X"d0",
X"bc",
X"4c",
X"3a",
X"f7",
X"a5",
X"fc",
X"d0",
X"0c",
X"a5",
X"fb",
X"d0",
X"2c",
X"ad",
X"b1",
X"07",
X"05",
X"f4",
X"d0",
X"ee",
X"60",
X"8d",
X"b1",
X"07",
X"c9",
X"01",
X"d0",
X"06",
X"20",
X"a7",
X"f4",
X"20",
X"71",
X"f5",
X"a6",
X"f4",
X"8e",
X"c5",
X"07",
X"a0",
X"00",
X"8c",
X"c4",
X"07",
X"84",
X"f4",
X"c9",
X"40",
X"d0",
X"30",
X"a2",
X"08",
X"8e",
X"c4",
X"07",
X"d0",
X"29",
X"c9",
X"04",
X"d0",
X"03",
X"20",
X"a7",
X"f4",
X"a0",
X"10",
X"8c",
X"c7",
X"07",
X"a0",
X"00",
X"8c",
X"b1",
X"07",
X"85",
X"f4",
X"c9",
X"01",
X"d0",
X"0e",
X"ee",
X"c7",
X"07",
X"ac",
X"c7",
X"07",
X"c0",
X"32",
X"d0",
X"0c",
X"a0",
X"11",
X"d0",
X"e4",
X"a0",
X"08",
X"84",
X"f7",
X"c8",
X"4a",
X"90",
X"fc",
X"b9",
X"0c",
X"f9",
X"a8",
X"b9",
X"0d",
X"f9",
X"85",
X"f0",
X"b9",
X"0e",
X"f9",
X"85",
X"f5",
X"b9",
X"0f",
X"f9",
X"85",
X"f6",
X"b9",
X"10",
X"f9",
X"85",
X"f9",
X"b9",
X"11",
X"f9",
X"85",
X"f8",
X"b9",
X"12",
X"f9",
X"8d",
X"b0",
X"07",
X"8d",
X"c1",
X"07",
X"a9",
X"01",
X"8d",
X"b4",
X"07",
X"8d",
X"b6",
X"07",
X"8d",
X"b9",
X"07",
X"8d",
X"ba",
X"07",
X"a9",
X"00",
X"85",
X"f7",
X"8d",
X"ca",
X"07",
X"a9",
X"0b",
X"8d",
X"15",
X"40",
X"a9",
X"0f",
X"8d",
X"15",
X"40",
X"ce",
X"b4",
X"07",
X"d0",
X"5f",
X"a4",
X"f7",
X"e6",
X"f7",
X"b1",
X"f5",
X"f0",
X"04",
X"10",
X"3d",
X"d0",
X"2f",
X"ad",
X"b1",
X"07",
X"c9",
X"40",
X"d0",
X"05",
X"ad",
X"c5",
X"07",
X"d0",
X"1d",
X"29",
X"04",
X"d0",
X"1c",
X"a5",
X"f4",
X"29",
X"5f",
X"d0",
X"13",
X"a9",
X"00",
X"85",
X"f4",
X"8d",
X"b1",
X"07",
X"8d",
X"08",
X"40",
X"a9",
X"90",
X"8d",
X"00",
X"40",
X"8d",
X"04",
X"40",
X"60",
X"4c",
X"d4",
X"f6",
X"4c",
X"a4",
X"f6",
X"20",
X"cb",
X"f8",
X"8d",
X"b3",
X"07",
X"a4",
X"f7",
X"e6",
X"f7",
X"b1",
X"f5",
X"a6",
X"f2",
X"d0",
X"0e",
X"20",
X"a9",
X"f3",
X"f0",
X"03",
X"20",
X"d8",
X"f8",
X"8d",
X"b5",
X"07",
X"20",
X"9f",
X"f3",
X"ad",
X"b3",
X"07",
X"8d",
X"b4",
X"07",
X"a5",
X"f2",
X"d0",
X"1a",
X"ad",
X"b1",
X"07",
X"29",
X"91",
X"d0",
X"13",
X"ac",
X"b5",
X"07",
X"f0",
X"03",
X"ce",
X"b5",
X"07",
X"20",
X"f4",
X"f8",
X"8d",
X"04",
X"40",
X"a2",
X"7f",
X"8e",
X"05",
X"40",
X"a4",
X"f8",
X"f0",
X"5a",
X"ce",
X"b6",
X"07",
X"d0",
X"32",
X"a4",
X"f8",
X"e6",
X"f8",
X"b1",
X"f5",
X"d0",
X"0f",
X"a9",
X"83",
X"8d",
X"00",
X"40",
X"a9",
X"94",
X"8d",
X"01",
X"40",
X"8d",
X"ca",
X"07",
X"d0",
X"e9",
X"20",
X"c5",
X"f8",
X"8d",
X"b6",
X"07",
X"a4",
X"f1",
X"d0",
X"34",
X"8a",
X"29",
X"3e",
X"20",
X"8b",
X"f3",
X"f0",
X"03",
X"20",
X"d8",
X"f8",
X"8d",
X"b7",
X"07",
X"20",
X"81",
X"f3",
X"a5",
X"f1",
X"d0",
X"1f",
X"ad",
X"b1",
X"07",
X"29",
X"91",
X"d0",
X"0e",
X"ac",
X"b7",
X"07",
X"f0",
X"03",
X"ce",
X"b7",
X"07",
X"20",
X"f4",
X"f8",
X"8d",
X"00",
X"40",
X"ad",
X"ca",
X"07",
X"d0",
X"02",
X"a9",
X"7f",
X"8d",
X"01",
X"40",
X"a5",
X"f9",
X"ce",
X"b9",
X"07",
X"d0",
X"4c",
X"a4",
X"f9",
X"e6",
X"f9",
X"b1",
X"f5",
X"f0",
X"41",
X"10",
X"13",
X"20",
X"cb",
X"f8",
X"8d",
X"b8",
X"07",
X"a9",
X"1f",
X"8d",
X"08",
X"40",
X"a4",
X"f9",
X"e6",
X"f9",
X"b1",
X"f5",
X"f0",
X"2c",
X"20",
X"ad",
X"f3",
X"ae",
X"b8",
X"07",
X"8e",
X"b9",
X"07",
X"ad",
X"b1",
X"07",
X"29",
X"6e",
X"d0",
X"06",
X"a5",
X"f4",
X"29",
X"0a",
X"f0",
X"19",
X"8a",
X"c9",
X"12",
X"b0",
X"0f",
X"ad",
X"b1",
X"07",
X"29",
X"08",
X"f0",
X"04",
X"a9",
X"0f",
X"d0",
X"06",
X"a9",
X"1f",
X"d0",
X"02",
X"a9",
X"ff",
X"8d",
X"08",
X"40",
X"a5",
X"f4",
X"29",
X"f3",
X"f0",
X"51",
X"ce",
X"ba",
X"07",
X"d0",
X"4c",
X"ac",
X"b0",
X"07",
X"ee",
X"b0",
X"07",
X"b1",
X"f5",
X"d0",
X"08",
X"ad",
X"c1",
X"07",
X"8d",
X"b0",
X"07",
X"d0",
X"ee",
X"20",
X"c5",
X"f8",
X"8d",
X"ba",
X"07",
X"8a",
X"29",
X"3e",
X"f0",
X"24",
X"c9",
X"30",
X"f0",
X"18",
X"c9",
X"20",
X"f0",
X"0c",
X"29",
X"10",
X"f0",
X"18",
X"a9",
X"1c",
X"a2",
X"03",
X"a0",
X"18",
X"d0",
X"12",
X"a9",
X"1c",
X"a2",
X"0c",
X"a0",
X"18",
X"d0",
X"0a",
X"a9",
X"1c",
X"a2",
X"03",
X"a0",
X"58",
X"d0",
X"02",
X"a9",
X"10",
X"8d",
X"0c",
X"40",
X"8e",
X"0e",
X"40",
X"8c",
X"0f",
X"40",
X"60",
X"aa",
X"6a",
X"8a",
X"2a",
X"2a",
X"2a",
X"29",
X"07",
X"18",
X"65",
X"f0",
X"6d",
X"c4",
X"07",
X"a8",
X"b9",
X"66",
X"ff",
X"60",
X"ad",
X"b1",
X"07",
X"29",
X"08",
X"f0",
X"04",
X"a9",
X"04",
X"d0",
X"0c",
X"a5",
X"f4",
X"29",
X"7d",
X"f0",
X"04",
X"a9",
X"08",
X"d0",
X"02",
X"a9",
X"28",
X"a2",
X"82",
X"a0",
X"7f",
X"60",
X"ad",
X"b1",
X"07",
X"29",
X"08",
X"f0",
X"04",
X"b9",
X"96",
X"ff",
X"60",
X"a5",
X"f4",
X"29",
X"7d",
X"f0",
X"04",
X"b9",
X"9a",
X"ff",
X"60",
X"b9",
X"a2",
X"ff",
X"60",
X"a5",
X"59",
X"54",
X"64",
X"59",
X"3c",
X"31",
X"4b",
X"69",
X"5e",
X"46",
X"4f",
X"36",
X"8d",
X"36",
X"4b",
X"8d",
X"69",
X"69",
X"6f",
X"75",
X"6f",
X"7b",
X"6f",
X"75",
X"6f",
X"7b",
X"81",
X"87",
X"81",
X"8d",
X"69",
X"69",
X"93",
X"99",
X"93",
X"9f",
X"93",
X"99",
X"93",
X"9f",
X"81",
X"87",
X"81",
X"8d",
X"93",
X"99",
X"93",
X"9f",
X"08",
X"72",
X"fc",
X"27",
X"18",
X"20",
X"b8",
X"f9",
X"2e",
X"1a",
X"40",
X"20",
X"b0",
X"fc",
X"3d",
X"21",
X"20",
X"c4",
X"fc",
X"3f",
X"1d",
X"18",
X"11",
X"fd",
X"00",
X"00",
X"08",
X"1c",
X"fa",
X"00",
X"00",
X"a4",
X"fb",
X"93",
X"62",
X"10",
X"c8",
X"fe",
X"24",
X"14",
X"18",
X"45",
X"fc",
X"1e",
X"14",
X"08",
X"52",
X"fd",
X"a0",
X"70",
X"68",
X"08",
X"51",
X"fe",
X"4c",
X"24",
X"18",
X"01",
X"fa",
X"2d",
X"1c",
X"b8",
X"18",
X"49",
X"fa",
X"20",
X"12",
X"70",
X"18",
X"75",
X"fa",
X"1b",
X"10",
X"44",
X"18",
X"9d",
X"fa",
X"11",
X"0a",
X"1c",
X"18",
X"c2",
X"fa",
X"2d",
X"10",
X"58",
X"18",
X"db",
X"fa",
X"14",
X"0d",
X"3f",
X"18",
X"f9",
X"fa",
X"15",
X"0d",
X"21",
X"18",
X"25",
X"fb",
X"18",
X"10",
X"7a",
X"18",
X"4b",
X"fb",
X"19",
X"0f",
X"54",
X"18",
X"74",
X"fb",
X"1e",
X"12",
X"2b",
X"18",
X"72",
X"fb",
X"1e",
X"0f",
X"2d",
X"84",
X"2c",
X"2c",
X"2c",
X"82",
X"04",
X"2c",
X"04",
X"85",
X"2c",
X"84",
X"2c",
X"2c",
X"2a",
X"2a",
X"2a",
X"82",
X"04",
X"2a",
X"04",
X"85",
X"2a",
X"84",
X"2a",
X"2a",
X"00",
X"1f",
X"1f",
X"1f",
X"98",
X"1f",
X"1f",
X"98",
X"9e",
X"98",
X"1f",
X"1d",
X"1d",
X"1d",
X"94",
X"1d",
X"1d",
X"94",
X"9c",
X"94",
X"1d",
X"86",
X"18",
X"85",
X"26",
X"30",
X"84",
X"04",
X"26",
X"30",
X"86",
X"14",
X"85",
X"22",
X"2c",
X"84",
X"04",
X"22",
X"2c",
X"21",
X"d0",
X"c4",
X"d0",
X"31",
X"d0",
X"c4",
X"d0",
X"00",
X"85",
X"2c",
X"22",
X"1c",
X"84",
X"26",
X"2a",
X"82",
X"28",
X"26",
X"04",
X"87",
X"22",
X"34",
X"3a",
X"82",
X"40",
X"04",
X"36",
X"84",
X"3a",
X"34",
X"82",
X"2c",
X"30",
X"85",
X"2a",
X"00",
X"5d",
X"55",
X"4d",
X"15",
X"19",
X"96",
X"15",
X"d5",
X"e3",
X"eb",
X"2d",
X"a6",
X"2b",
X"27",
X"9c",
X"9e",
X"59",
X"85",
X"22",
X"1c",
X"14",
X"84",
X"1e",
X"22",
X"82",
X"20",
X"1e",
X"04",
X"87",
X"1c",
X"2c",
X"34",
X"82",
X"36",
X"04",
X"30",
X"34",
X"04",
X"2c",
X"04",
X"26",
X"2a",
X"85",
X"22",
X"84",
X"04",
X"82",
X"3a",
X"38",
X"36",
X"32",
X"04",
X"34",
X"04",
X"24",
X"26",
X"2c",
X"04",
X"26",
X"2c",
X"30",
X"00",
X"05",
X"b4",
X"b2",
X"b0",
X"2b",
X"ac",
X"84",
X"9c",
X"9e",
X"a2",
X"84",
X"94",
X"9c",
X"9e",
X"85",
X"14",
X"22",
X"84",
X"2c",
X"85",
X"1e",
X"82",
X"2c",
X"84",
X"2c",
X"1e",
X"84",
X"04",
X"82",
X"3a",
X"38",
X"36",
X"32",
X"04",
X"34",
X"04",
X"64",
X"04",
X"64",
X"86",
X"64",
X"00",
X"05",
X"b4",
X"b2",
X"b0",
X"2b",
X"ac",
X"84",
X"37",
X"b6",
X"b6",
X"45",
X"85",
X"14",
X"1c",
X"82",
X"22",
X"84",
X"2c",
X"4e",
X"82",
X"4e",
X"84",
X"4e",
X"22",
X"84",
X"04",
X"85",
X"32",
X"85",
X"30",
X"86",
X"2c",
X"04",
X"00",
X"05",
X"a4",
X"05",
X"9e",
X"05",
X"9d",
X"85",
X"84",
X"14",
X"85",
X"24",
X"28",
X"2c",
X"82",
X"22",
X"84",
X"22",
X"14",
X"21",
X"d0",
X"c4",
X"d0",
X"31",
X"d0",
X"c4",
X"d0",
X"00",
X"82",
X"2c",
X"84",
X"2c",
X"2c",
X"82",
X"2c",
X"30",
X"04",
X"34",
X"2c",
X"04",
X"26",
X"86",
X"22",
X"00",
X"a4",
X"25",
X"25",
X"a4",
X"29",
X"a2",
X"1d",
X"9c",
X"95",
X"82",
X"2c",
X"2c",
X"04",
X"2c",
X"04",
X"2c",
X"30",
X"85",
X"34",
X"04",
X"04",
X"00",
X"a4",
X"25",
X"25",
X"a4",
X"a8",
X"63",
X"04",
X"85",
X"0e",
X"1a",
X"84",
X"24",
X"85",
X"22",
X"14",
X"84",
X"0c",
X"82",
X"34",
X"84",
X"34",
X"34",
X"82",
X"2c",
X"84",
X"34",
X"86",
X"3a",
X"04",
X"00",
X"a0",
X"21",
X"21",
X"a0",
X"21",
X"2b",
X"05",
X"a3",
X"82",
X"18",
X"84",
X"18",
X"18",
X"82",
X"18",
X"18",
X"04",
X"86",
X"3a",
X"22",
X"31",
X"90",
X"31",
X"90",
X"31",
X"71",
X"31",
X"90",
X"90",
X"90",
X"00",
X"82",
X"34",
X"84",
X"2c",
X"85",
X"22",
X"84",
X"24",
X"82",
X"26",
X"36",
X"04",
X"36",
X"86",
X"26",
X"00",
X"ac",
X"27",
X"5d",
X"1d",
X"9e",
X"2d",
X"ac",
X"9f",
X"85",
X"14",
X"82",
X"20",
X"84",
X"22",
X"2c",
X"1e",
X"1e",
X"82",
X"2c",
X"2c",
X"1e",
X"04",
X"87",
X"2a",
X"40",
X"40",
X"40",
X"3a",
X"36",
X"82",
X"34",
X"2c",
X"04",
X"26",
X"86",
X"22",
X"00",
X"e3",
X"f7",
X"f7",
X"f7",
X"f5",
X"f1",
X"ac",
X"27",
X"9e",
X"9d",
X"85",
X"18",
X"82",
X"1e",
X"84",
X"22",
X"2a",
X"22",
X"22",
X"82",
X"2c",
X"2c",
X"22",
X"04",
X"86",
X"04",
X"82",
X"2a",
X"36",
X"04",
X"36",
X"87",
X"36",
X"34",
X"30",
X"86",
X"2c",
X"04",
X"00",
X"00",
X"68",
X"6a",
X"6c",
X"45",
X"a2",
X"31",
X"b0",
X"f1",
X"ed",
X"eb",
X"a2",
X"1d",
X"9c",
X"95",
X"86",
X"04",
X"85",
X"22",
X"82",
X"22",
X"87",
X"22",
X"26",
X"2a",
X"84",
X"2c",
X"22",
X"86",
X"14",
X"51",
X"90",
X"31",
X"11",
X"00",
X"80",
X"22",
X"28",
X"22",
X"26",
X"22",
X"24",
X"22",
X"26",
X"22",
X"28",
X"22",
X"2a",
X"22",
X"28",
X"22",
X"26",
X"22",
X"28",
X"22",
X"26",
X"22",
X"24",
X"22",
X"26",
X"22",
X"28",
X"22",
X"2a",
X"22",
X"28",
X"22",
X"26",
X"20",
X"26",
X"20",
X"24",
X"20",
X"26",
X"20",
X"28",
X"20",
X"26",
X"20",
X"28",
X"20",
X"26",
X"20",
X"24",
X"20",
X"26",
X"20",
X"24",
X"20",
X"26",
X"20",
X"28",
X"20",
X"26",
X"20",
X"28",
X"20",
X"26",
X"20",
X"24",
X"28",
X"30",
X"28",
X"32",
X"28",
X"30",
X"28",
X"2e",
X"28",
X"30",
X"28",
X"2e",
X"28",
X"2c",
X"28",
X"2e",
X"28",
X"30",
X"28",
X"32",
X"28",
X"30",
X"28",
X"2e",
X"28",
X"30",
X"28",
X"2e",
X"28",
X"2c",
X"28",
X"2e",
X"00",
X"04",
X"70",
X"6e",
X"6c",
X"6e",
X"70",
X"72",
X"70",
X"6e",
X"70",
X"6e",
X"6c",
X"6e",
X"70",
X"72",
X"70",
X"6e",
X"6e",
X"6c",
X"6e",
X"70",
X"6e",
X"70",
X"6e",
X"6c",
X"6e",
X"6c",
X"6e",
X"70",
X"6e",
X"70",
X"6e",
X"6c",
X"76",
X"78",
X"76",
X"74",
X"76",
X"74",
X"72",
X"74",
X"76",
X"78",
X"76",
X"74",
X"76",
X"74",
X"72",
X"74",
X"84",
X"1a",
X"83",
X"18",
X"20",
X"84",
X"1e",
X"83",
X"1c",
X"28",
X"26",
X"1c",
X"1a",
X"1c",
X"82",
X"2c",
X"04",
X"04",
X"22",
X"04",
X"04",
X"84",
X"1c",
X"87",
X"26",
X"2a",
X"26",
X"84",
X"24",
X"28",
X"24",
X"80",
X"22",
X"00",
X"9c",
X"05",
X"94",
X"05",
X"0d",
X"9f",
X"1e",
X"9c",
X"98",
X"9d",
X"82",
X"22",
X"04",
X"04",
X"1c",
X"04",
X"04",
X"84",
X"14",
X"86",
X"1e",
X"80",
X"16",
X"80",
X"14",
X"81",
X"1c",
X"30",
X"04",
X"30",
X"30",
X"04",
X"1e",
X"32",
X"04",
X"32",
X"32",
X"04",
X"20",
X"34",
X"04",
X"34",
X"34",
X"04",
X"36",
X"04",
X"84",
X"36",
X"00",
X"46",
X"a4",
X"64",
X"a4",
X"48",
X"a6",
X"66",
X"a6",
X"4a",
X"a8",
X"68",
X"a8",
X"6a",
X"44",
X"2b",
X"81",
X"2a",
X"42",
X"04",
X"42",
X"42",
X"04",
X"2c",
X"64",
X"04",
X"64",
X"64",
X"04",
X"2e",
X"46",
X"04",
X"46",
X"46",
X"04",
X"22",
X"04",
X"84",
X"22",
X"87",
X"04",
X"06",
X"0c",
X"14",
X"1c",
X"22",
X"86",
X"2c",
X"22",
X"87",
X"04",
X"60",
X"0e",
X"14",
X"1a",
X"24",
X"86",
X"2c",
X"24",
X"87",
X"04",
X"08",
X"10",
X"18",
X"1e",
X"28",
X"86",
X"30",
X"30",
X"80",
X"64",
X"00",
X"cd",
X"d5",
X"dd",
X"e3",
X"ed",
X"f5",
X"bb",
X"b5",
X"cf",
X"d5",
X"db",
X"e5",
X"ed",
X"f3",
X"bd",
X"b3",
X"d1",
X"d9",
X"df",
X"e9",
X"f1",
X"f7",
X"bf",
X"ff",
X"ff",
X"ff",
X"34",
X"00",
X"86",
X"04",
X"87",
X"14",
X"1c",
X"22",
X"86",
X"34",
X"84",
X"2c",
X"04",
X"04",
X"04",
X"87",
X"14",
X"1a",
X"24",
X"86",
X"32",
X"84",
X"2c",
X"04",
X"86",
X"04",
X"87",
X"18",
X"1e",
X"28",
X"86",
X"36",
X"87",
X"30",
X"30",
X"30",
X"80",
X"2c",
X"82",
X"14",
X"2c",
X"62",
X"26",
X"10",
X"28",
X"80",
X"04",
X"82",
X"14",
X"2c",
X"62",
X"26",
X"10",
X"28",
X"80",
X"04",
X"82",
X"08",
X"1e",
X"5e",
X"18",
X"60",
X"1a",
X"80",
X"04",
X"82",
X"08",
X"1e",
X"5e",
X"18",
X"60",
X"1a",
X"86",
X"04",
X"83",
X"1a",
X"18",
X"16",
X"84",
X"14",
X"1a",
X"18",
X"0e",
X"0c",
X"16",
X"83",
X"14",
X"20",
X"1e",
X"1c",
X"28",
X"26",
X"87",
X"24",
X"1a",
X"12",
X"10",
X"62",
X"0e",
X"80",
X"04",
X"04",
X"00",
X"82",
X"18",
X"1c",
X"20",
X"22",
X"26",
X"28",
X"81",
X"2a",
X"2a",
X"2a",
X"04",
X"2a",
X"04",
X"83",
X"2a",
X"82",
X"22",
X"86",
X"34",
X"32",
X"34",
X"81",
X"04",
X"22",
X"26",
X"2a",
X"2c",
X"30",
X"86",
X"34",
X"83",
X"32",
X"82",
X"36",
X"84",
X"34",
X"85",
X"04",
X"81",
X"22",
X"86",
X"30",
X"2e",
X"30",
X"81",
X"04",
X"22",
X"26",
X"2a",
X"2c",
X"2e",
X"86",
X"30",
X"83",
X"22",
X"82",
X"36",
X"84",
X"34",
X"85",
X"04",
X"81",
X"22",
X"86",
X"3a",
X"3a",
X"3a",
X"82",
X"3a",
X"81",
X"40",
X"82",
X"04",
X"81",
X"3a",
X"86",
X"36",
X"36",
X"36",
X"82",
X"36",
X"81",
X"3a",
X"82",
X"04",
X"81",
X"36",
X"86",
X"34",
X"82",
X"26",
X"2a",
X"36",
X"81",
X"34",
X"34",
X"85",
X"34",
X"81",
X"2a",
X"86",
X"2c",
X"00",
X"84",
X"90",
X"b0",
X"84",
X"50",
X"50",
X"b0",
X"00",
X"98",
X"96",
X"94",
X"92",
X"94",
X"96",
X"58",
X"58",
X"58",
X"44",
X"5c",
X"44",
X"9f",
X"a3",
X"a1",
X"a3",
X"85",
X"a3",
X"e0",
X"a6",
X"23",
X"c4",
X"9f",
X"9d",
X"9f",
X"85",
X"9f",
X"d2",
X"a6",
X"23",
X"c4",
X"b5",
X"b1",
X"af",
X"85",
X"b1",
X"af",
X"ad",
X"85",
X"95",
X"9e",
X"a2",
X"aa",
X"6a",
X"6a",
X"6b",
X"5e",
X"9d",
X"84",
X"04",
X"04",
X"82",
X"22",
X"86",
X"22",
X"82",
X"14",
X"22",
X"2c",
X"12",
X"22",
X"2a",
X"14",
X"22",
X"2c",
X"1c",
X"22",
X"2c",
X"14",
X"22",
X"2c",
X"12",
X"22",
X"2a",
X"14",
X"22",
X"2c",
X"1c",
X"22",
X"2c",
X"18",
X"22",
X"2a",
X"16",
X"20",
X"28",
X"18",
X"22",
X"2a",
X"12",
X"22",
X"2a",
X"18",
X"22",
X"2a",
X"12",
X"22",
X"2a",
X"14",
X"22",
X"2c",
X"0c",
X"22",
X"2c",
X"14",
X"22",
X"34",
X"12",
X"22",
X"30",
X"10",
X"22",
X"2e",
X"16",
X"22",
X"34",
X"18",
X"26",
X"36",
X"16",
X"26",
X"36",
X"14",
X"26",
X"36",
X"12",
X"22",
X"36",
X"5c",
X"22",
X"34",
X"0c",
X"22",
X"22",
X"81",
X"1e",
X"1e",
X"85",
X"1e",
X"81",
X"12",
X"86",
X"14",
X"81",
X"2c",
X"22",
X"1c",
X"2c",
X"22",
X"1c",
X"85",
X"2c",
X"04",
X"81",
X"2e",
X"24",
X"1e",
X"2e",
X"24",
X"1e",
X"85",
X"2e",
X"04",
X"81",
X"32",
X"28",
X"22",
X"32",
X"28",
X"22",
X"85",
X"32",
X"87",
X"36",
X"36",
X"36",
X"84",
X"3a",
X"00",
X"5c",
X"54",
X"4c",
X"5c",
X"54",
X"4c",
X"5c",
X"1c",
X"1c",
X"5c",
X"5c",
X"5c",
X"5c",
X"5e",
X"56",
X"4e",
X"5e",
X"56",
X"4e",
X"5e",
X"1e",
X"1e",
X"5e",
X"5e",
X"5e",
X"5e",
X"62",
X"5a",
X"50",
X"62",
X"5a",
X"50",
X"62",
X"22",
X"22",
X"62",
X"e7",
X"e7",
X"e7",
X"2b",
X"86",
X"14",
X"81",
X"14",
X"80",
X"14",
X"14",
X"81",
X"14",
X"14",
X"14",
X"14",
X"86",
X"16",
X"81",
X"16",
X"80",
X"16",
X"16",
X"81",
X"16",
X"16",
X"16",
X"16",
X"81",
X"28",
X"22",
X"1a",
X"28",
X"22",
X"1a",
X"28",
X"80",
X"28",
X"28",
X"81",
X"28",
X"87",
X"2c",
X"2c",
X"2c",
X"84",
X"30",
X"83",
X"04",
X"84",
X"0c",
X"83",
X"62",
X"10",
X"84",
X"12",
X"83",
X"1c",
X"22",
X"1e",
X"22",
X"26",
X"18",
X"1e",
X"04",
X"1c",
X"00",
X"e3",
X"e1",
X"e3",
X"1d",
X"de",
X"e0",
X"23",
X"ec",
X"75",
X"74",
X"f0",
X"f4",
X"f6",
X"ea",
X"31",
X"2d",
X"83",
X"12",
X"14",
X"04",
X"18",
X"1a",
X"1c",
X"14",
X"26",
X"22",
X"1e",
X"1c",
X"18",
X"1e",
X"22",
X"0c",
X"14",
X"ff",
X"ff",
X"ff",
X"00",
X"88",
X"00",
X"2f",
X"00",
X"00",
X"02",
X"a6",
X"02",
X"80",
X"02",
X"5c",
X"02",
X"3a",
X"02",
X"1a",
X"01",
X"df",
X"01",
X"c4",
X"01",
X"ab",
X"01",
X"93",
X"01",
X"7c",
X"01",
X"67",
X"01",
X"53",
X"01",
X"40",
X"01",
X"2e",
X"01",
X"1d",
X"01",
X"0d",
X"00",
X"fe",
X"00",
X"ef",
X"00",
X"e2",
X"00",
X"d5",
X"00",
X"c9",
X"00",
X"be",
X"00",
X"b3",
X"00",
X"a9",
X"00",
X"a0",
X"00",
X"97",
X"00",
X"8e",
X"00",
X"86",
X"00",
X"77",
X"00",
X"7e",
X"00",
X"71",
X"00",
X"54",
X"00",
X"64",
X"00",
X"5f",
X"00",
X"59",
X"00",
X"50",
X"00",
X"47",
X"00",
X"43",
X"00",
X"3b",
X"00",
X"35",
X"00",
X"2a",
X"00",
X"23",
X"04",
X"75",
X"03",
X"57",
X"02",
X"f9",
X"02",
X"cf",
X"01",
X"fc",
X"00",
X"6a",
X"05",
X"0a",
X"14",
X"28",
X"50",
X"1e",
X"3c",
X"02",
X"04",
X"08",
X"10",
X"20",
X"40",
X"18",
X"30",
X"0c",
X"03",
X"06",
X"0c",
X"18",
X"30",
X"12",
X"24",
X"08",
X"36",
X"03",
X"09",
X"06",
X"12",
X"1b",
X"24",
X"0c",
X"24",
X"02",
X"06",
X"04",
X"0c",
X"12",
X"18",
X"08",
X"12",
X"01",
X"03",
X"02",
X"06",
X"09",
X"0c",
X"04",
X"98",
X"99",
X"9a",
X"9b",
X"90",
X"94",
X"94",
X"95",
X"95",
X"96",
X"97",
X"98",
X"90",
X"91",
X"92",
X"92",
X"93",
X"93",
X"93",
X"94",
X"94",
X"94",
X"94",
X"94",
X"94",
X"95",
X"95",
X"95",
X"95",
X"95",
X"95",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"96",
X"95",
X"95",
X"94",
X"93",
X"15",
X"16",
X"16",
X"17",
X"17",
X"18",
X"19",
X"19",
X"1a",
X"1a",
X"1c",
X"1d",
X"1d",
X"1e",
X"1e",
X"1f",
X"1f",
X"1f",
X"1f",
X"1e",
X"1d",
X"1c",
X"1e",
X"1f",
X"1f",
X"1e",
X"1d",
X"1c",
X"1a",
X"18",
X"16",
X"14",
X"15",
X"16",
X"16",
X"17",
X"17",
X"18",
X"19",
X"19",
X"1a",
X"1a",
X"1c",
X"1d",
X"1d",
X"1e",
X"1e",
X"1f",
X"82",
X"80",
X"00",
X"80",
X"f0",
X"ff"
);
	
begin
	
	process(clock)
	begin
		if(rising_edge(clock)) then
			q <= rom(address);
		end if;
	end process;
		
end rtl;
